library ieee ;
    use ieee.std_logic_1164.all ;
    use ieee.numeric_std.all ;
    use IEEE.std_logic_arith.all;
    use IEEE.std_logic_unsigned.all;

entity UC is
    generic (
        wl_Q:   integer:= 4;
        wl_T:   integer:= 4
    );
  port (
    q_in:   in  std_logic_vector(wl_Q-1 downto 0);
    t_in:   in  std_logic_vector(wl_T-1 downto 0);
    c_in:   in  std_logic;
  --  z_in:   in  std_logic;
    Xs_out: out std_logic_vector(9 downto 0)
    --x0, x1, x2, x3, x4, x5, x6, x7, x8, x9: out std_logic
  ) ;
end UC ; 
--:= (others => '0' )
architecture arch of UC is

    signal control : std_logic_vector(7 downto 0);  -- control de entradas
    signal  x0, x1, x2, x3, x5, x6, x7, x8, x9:  std_logic;
    --signal xs: std_logic_vector(wl_Xs downto 0); -- array salida xs
    --signal flags: std_logic_vector(1 downto 0);-- entradas banderas
begin
    
   control <= q_in & t_in; -- concatenando entradas q y t

    process (q_in, t_in, control )
    begin
        case( control ) is
------------  00h  MOV A, N
        --       q & t
            when "00000000" => --t0
                x0  <= '0';
                x1  <= '0';
                x2  <= '0';
                x3  <= '0';
                x5  <= '0';
                x6  <= '0';
                x7  <= '0';
                x8  <= '1';
                x9  <= '0';


            when "00000001" => --t1
                x0  <= '0';
                x1  <= '0';
                x2  <= '1';
                x3  <= '0';
                x5  <= '0';
                x6  <= '1';
                x7  <= '0';
                x8  <= '0';
                x9  <= '0';
    
                
            when "00000010" => --t2
                x0  <= '1';
                x1  <= '0';
                x2  <= '0';
                x3  <= '0';
                x5  <= '0';
                x6  <= '0';
                x7  <= '0';
                x8  <= '0';
                x9  <= '0';
    
                
            when "00000011" => --t3q0
                x0  <= '0';
                x1  <= '0';
                x2  <= '0';
                x3  <= '0';
                x5  <= '0';
                x6  <= '0';
                x7  <= '0';
                x8  <= '1';
                x9  <= '0';
  
                
            when "00000100" => --t4q0
                x0  <= '0';
                x1  <= '0';
                x2  <= '1';
                x3  <= '0';
                x5  <= '0';
                x6  <= '1';
                x7  <= '0';
                x8  <= '0';
                x9  <= '0';
   

            when "00000101" => --t5q0
                x0  <= '0';
                x1  <= '0';
                x2  <= '0';
                x3  <= '0';
                x5  <= '0';
                x6  <= '0';
                x7  <= '0';
                x8  <= '0';
                x9  <= '0';
 
            
            when "00000110" => --t6q0
                x0  <= '0';
                x1  <= '0';
                x2  <= '0';
                x3  <= '0';
                x5  <= '0';
                x6  <= '0';
                x7  <= '0';
                x8  <= '0';
                x9  <= '0';
         
------------  FIN -> 00h  MOV A, N            
            
------------  01h  MOV A, [DIR]
        --       q & t
            when "00010000" => --t0
                x0  <= '0';
                x1  <= '0';
                x2  <= '0';
                x3  <= '0';
                x5  <= '0';
                x6  <= '0';
                x7  <= '0';
                x8  <= '1';
                x9  <= '0';


            when "00010001" => --t1
                x0  <= '0';
                x1  <= '0';
                x2  <= '1';
                x3  <= '0';
                x5  <= '0';
                x6  <= '1';
                x7  <= '0';
                x8  <= '0';
                x9  <= '0';
    

            when "00010010" => --t2
                x0  <= '1';
                x1  <= '0';
                x2  <= '0';
                x3  <= '0';
                x5  <= '0';
                x6  <= '0';
                x7  <= '0';
                x8  <= '0';
                x9  <= '0';
    

            when "00010011" => --t3q1
                x0  <= '0';
                x1  <= '0';
                x2  <= '0';
                x3  <= '0';
                x5  <= '0';
                x6  <= '0';
                x7  <= '0';
                x8  <= '1';
                x9  <= '0';
  

            when "00010100" => --t4q1
                x0  <= '0';
                x1  <= '0';
                x2  <= '1';
                x3  <= '0';
                x5  <= '0';
                x6  <= '1';
                x7  <= '0';
                x8  <= '0';
                x9  <= '0';
   

            when "00010101" => --t5q1
                x0  <= '0';
                x1  <= '0';
                x2  <= '0';
                x3  <= '0';
                x5  <= '0';
                x6  <= '0';
                x7  <= '0';
                x8  <= '0';
                x9  <= '0';
 

            when "00010110" => --t6q1
                x0  <= '0';
                x1  <= '0';
                x2  <= '0';
                x3  <= '0';
                x5  <= '0';
                x6  <= '0';
                x7  <= '0';
                x8  <= '1';
                x9  <= '0';

                
            when "00010111" => --t7q1
                x0  <= '0';
                x1  <= '0';
                x2  <= '1';
                x3  <= '0';
                x5  <= '0';
                x6  <= '1';
                x7  <= '0';
                x8  <= '0';
                x9  <= '0';

                
            when "00011000" => --t8q1
                x0  <= '0';
                x1  <= '0';
                x2  <= '0';
                x3  <= '0';
                x5  <= '0';
                x6  <= '0';
                x7  <= '1';
                x8  <= '0';
                x9  <= '0';

                
            when "00011001" => --t9q1
                x0  <= '0';
                x1  <= '0';
                x2  <= '1';
                x3  <= '0';
                x5  <= '0';
                x6  <= '0';
                x7  <= '0';
                x8  <= '0';
                x9  <= '0';

            when "00011010" => --tAq1 
                x0  <= '0';
                x1  <= '0';
                x2  <= '0';
                x3  <= '0';
                x5  <= '0';
                x6  <= '0';
                x7  <= '0';
                x8  <= '0';
                x9  <= '0';


            when "00011011" => --tBq1
                x0  <= '0';
                x1  <= '0';
                x2  <= '0';
                x3  <= '0';
                x5  <= '0';
                x6  <= '0';
                x7  <= '0';
                x8  <= '0';
                x9  <= '0';


------------  FIN -> MOV A, [DIR]           
    
------------ 02h  MOV SP, [N]
        --       q & t
        when "00100000" => --t0
            x0  <= '0';
            x1  <= '0';
            x2  <= '0';
            x3  <= '0';
            x5  <= '0';
            x6  <= '0';
            x7  <= '0';
            x8  <= '1';
            x9  <= '0';

        when "00100001" => --t1
            x0  <= '0';
            x1  <= '0';
            x2  <= '1';
            x3  <= '0';
            x5  <= '0';
            x6  <= '1';
            x7  <= '0';
            x8  <= '0';
            x9  <= '0';    
            
        when "00100010" => --t2
            x0  <= '1';
            x1  <= '0';
            x2  <= '0';
            x3  <= '0';
            x5  <= '0';
            x6  <= '0';
            x7  <= '0';
            x8  <= '0';
            x9  <= '0';    
            
        when "00100011" => --t3q2
            x0  <= '0';
            x1  <= '0';
            x2  <= '0';
            x3  <= '0';
            x5  <= '0';
            x6  <= '0';
            x7  <= '0';
            x8  <= '1';
            x9  <= '0';  
            
        when "00100100" => --t4q2
            x0  <= '0';
            x1  <= '0';
            x2  <= '1';
            x3  <= '0';
            x5  <= '0';
            x6  <= '1';
            x7  <= '0';
            x8  <= '0';
            x9  <= '0';   

        when "00100101" => --t5q2
            x0  <= '0';
            x1  <= '0';
            x2  <= '0';
            x3  <= '0';
            x5  <= '0';
            x6  <= '0';
            x7  <= '0';
            x8  <= '0';
            x9  <= '0'; 
            
        when "00100110" => --t6q2
            x0  <= '0';
            x1  <= '0';
            x2  <= '0';
            x3  <= '0';
            x5  <= '0';
            x6  <= '0';
            x7  <= '0';
            x8  <= '0';
            x9  <= '0';         
------------  FIN -> 02h  MOV SP, [N]           
            
------------ 03h  MOV [DIR], A
        --       q & t
        when "00110000" => --t0
            x0  <= '0';
            x1  <= '0';
            x2  <= '0';
            x3  <= '0';
            x5  <= '0';
            x6  <= '0';
            x7  <= '0';
            x8  <= '1';
            x9  <= '0';

        when "00110001" => --t1
            x0  <= '0';
            x1  <= '0';
            x2  <= '1';
            x3  <= '0';
            x5  <= '0';
            x6  <= '1';
            x7  <= '0';
            x8  <= '0';
            x9  <= '0';    
            
        when "00110010" => --t2
            x0  <= '1';
            x1  <= '0';
            x2  <= '0';
            x3  <= '0';
            x5  <= '0';
            x6  <= '0';
            x7  <= '0';
            x8  <= '0';
            x9  <= '0';    
            
        when "00110011" => --t3q3
            x0  <= '0';
            x1  <= '0';
            x2  <= '0';
            x3  <= '0';
            x5  <= '0';
            x6  <= '0';
            x7  <= '0';
            x8  <= '1';
            x9  <= '0';  
            
        when "00110100" => --t4q3
            x0  <= '0';
            x1  <= '0';
            x2  <= '1';
            x3  <= '0';
            x5  <= '0';
            x6  <= '1';
            x7  <= '0';
            x8  <= '0';
            x9  <= '0';   

        when "00110101" => --t5q3
            x0  <= '0';
            x1  <= '0';
            x2  <= '0';
            x3  <= '0';
            x5  <= '0';
            x6  <= '0';
            x7  <= '0';
            x8  <= '0';
            x9  <= '0'; 
            
        when "00110110" => --t6q3
            x0  <= '0';
            x1  <= '0';
            x2  <= '0';
            x3  <= '0';
            x5  <= '0';
            x6  <= '0';
            x7  <= '0';
            x8  <= '1';
            x9  <= '0'; 
            
        when "00110111" => --t7q3
            x0  <= '0';
            x1  <= '0';
            x2  <= '1';
            x3  <= '0';
            x5  <= '0';
            x6  <= '1';
            x7  <= '0';
            x8  <= '0';
            x9  <= '0'; 

        when "00111000" => --t8q3
            x0  <= '0';
            x1  <= '0';
            x2  <= '0';
            x3  <= '0';
            x5  <= '0';
            x6  <= '0';
            x7  <= '1';
            x8  <= '0';
            x9  <= '0'; 

        when "00111001" => --t9q3
            x0  <= '0';
            x1  <= '1';
            x2  <= '0';
            x3  <= '0';
            x5  <= '0';
            x6  <= '0';
            x7  <= '0';
            x8  <= '0';
            x9  <= '0'; 

        when "00111010" => --tAq3
            x0  <= '0';
            x1  <= '0';
            x2  <= '0';
            x3  <= '0';
            x5  <= '0';
            x6  <= '0';
            x7  <= '0';
            x8  <= '0';
            x9  <= '0'; 

        when "00111011" => --tBq3
            x0  <= '0';
            x1  <= '0';
            x2  <= '0';
            x3  <= '0';
            x5  <= '0';
            x6  <= '0';
            x7  <= '0';
            x8  <= '0';
            x9  <= '0'; 
------------  FIN -> 03h  MOV [DIR], A            
            
------------ 04h  XOR A, N     
        --       q & t
        when "01000000" => --t0
            x0  <= '0';
            x1  <= '0';
            x2  <= '0';
            x3  <= '0';
            x5  <= '0';
            x6  <= '0';
            x7  <= '0';
            x8  <= '1';
            x9  <= '0';

        when "01000001" => --t1
            x0  <= '0';
            x1  <= '0';
            x2  <= '1';
            x3  <= '0';
            x5  <= '0';
            x6  <= '1';
            x7  <= '0';
            x8  <= '0';
            x9  <= '0';    
            
        when "01000010" => --t2
            x0  <= '1';
            x1  <= '0';
            x2  <= '0';
            x3  <= '0';
            x5  <= '0';
            x6  <= '0';
            x7  <= '0';
            x8  <= '0';
            x9  <= '0';    
            
        when "01000011" => --t3q4
            x0  <= '0';
            x1  <= '0';
            x2  <= '0';
            x3  <= '0';
            x5  <= '0';
            x6  <= '0';
            x7  <= '0';
            x8  <= '1';
            x9  <= '0';  
            
        when "01000100" => --t4q4
            x0  <= '0';
            x1  <= '0';
            x2  <= '1';
            x3  <= '0';
            x5  <= '0';
            x6  <= '1';
            x7  <= '0';
            x8  <= '0';
            x9  <= '0';   

        when "01000101" => --t5q4
            x0  <= '0';
            x1  <= '0';
            x2  <= '0';
            x3  <= '0';
            x5  <= '0';
            x6  <= '0';
            x7  <= '0';
            x8  <= '0';
            x9  <= '0'; 
            
        when "01000110" => --t6q4
            x0  <= '0';
            x1  <= '0';
            x2  <= '0';
            x3  <= '0';
            x5  <= '0';
            x6  <= '0';
            x7  <= '0';
            x8  <= '0';
            x9  <= '0'; 
------------  FIN -> 04h  XOR A, N        
            
------------ 05h  ADD A, [DIR]    
        --       q & t
        when "01010000" => --t0
            x0  <= '0';
            x1  <= '0';
            x2  <= '0';
            x3  <= '0';
            x5  <= '0';
            x6  <= '0';
            x7  <= '0';
            x8  <= '1';
            x9  <= '0';

        when "01010001" => --t1
            x0  <= '0';
            x1  <= '0';
            x2  <= '1';
            x3  <= '0';
            x5  <= '0';
            x6  <= '1';
            x7  <= '0';
            x8  <= '0';
            x9  <= '0';    
            
        when "01010010" => --t2
            x0  <= '1';
            x1  <= '0';
            x2  <= '0';
            x3  <= '0';
            x5  <= '0';
            x6  <= '0';
            x7  <= '0';
            x8  <= '0';
            x9  <= '0';    
            
        when "01010011" => --t3q5
            x0  <= '0';
            x1  <= '0';
            x2  <= '0';
            x3  <= '0';
            x5  <= '0';
            x6  <= '0';
            x7  <= '0';
            x8  <= '1';
            x9  <= '0';  
            
        when "01010100" => --t4q5
            x0  <= '0';
            x1  <= '0';
            x2  <= '1';
            x3  <= '0';
            x5  <= '0';
            x6  <= '1';
            x7  <= '0';
            x8  <= '0';
            x9  <= '0';   

        when "01010101" => --t5q5
            x0  <= '0';
            x1  <= '0';
            x2  <= '0';
            x3  <= '0';
            x5  <= '0';
            x6  <= '0';
            x7  <= '0';
            x8  <= '0';
            x9  <= '0'; 
            
        when "01010110" => --t6q5
            x0  <= '0';
            x1  <= '0';
            x2  <= '0';
            x3  <= '0';
            x5  <= '0';
            x6  <= '0';
            x7  <= '0';
            x8  <= '1';
            x9  <= '0'; 

        when "01010111" => --t7q5
            x0  <= '0';
            x1  <= '0';
            x2  <= '1';
            x3  <= '0';
            x5  <= '0';
            x6  <= '1';
            x7  <= '0';
            x8  <= '0';
            x9  <= '0'; 

        when "01011000" => --t8q5
            x0  <= '0';
            x1  <= '0';
            x2  <= '0';
            x3  <= '0';
            x5  <= '0';
            x6  <= '0';
            x7  <= '1';
            x8  <= '0';
            x9  <= '0'; 

        when "01011001" => --t9q5
            x0  <= '0';
            x1  <= '0';
            x2  <= '1';
            x3  <= '0';
            x5  <= '0';
            x6  <= '0';
            x7  <= '0';
            x8  <= '0';
            x9  <= '0'; 

        when "01011010" => --tAq5
            x0  <= '0';
            x1  <= '0';
            x2  <= '0';
            x3  <= '0';
            x5  <= '0';
            x6  <= '0';
            x7  <= '0';
            x8  <= '0';
            x9  <= '0'; 

        when "01011011" => --tBq5
            x0  <= '0';
            x1  <= '0';
            x2  <= '0';
            x3  <= '0';
            x5  <= '0';
            x6  <= '0';
            x7  <= '0';
            x8  <= '0';
            x9  <= '0'; 
------------  FIN -> 05h  ADD A, [DIR]   
    
------------ 06h  AND A, [DIR]    
        --       q & t
        when "01100000" => --t0
            x0  <= '0';
            x1  <= '0';
            x2  <= '0';
            x3  <= '0';
            x5  <= '0';
            x6  <= '0';
            x7  <= '0';
            x8  <= '1';
            x9  <= '0';

        when "01100001" => --t1
            x0  <= '0';
            x1  <= '0';
            x2  <= '1';
            x3  <= '0';
            x5  <= '0';
            x6  <= '1';
            x7  <= '0';
            x8  <= '0';
            x9  <= '0';    
            
        when "01100010" => --t2
            x0  <= '1';
            x1  <= '0';
            x2  <= '0';
            x3  <= '0';
            x5  <= '0';
            x6  <= '0';
            x7  <= '0';
            x8  <= '0';
            x9  <= '0';    
            
        when "01100011" => --t3q6
            x0  <= '0';
            x1  <= '0';
            x2  <= '1';
            x3  <= '0';
            x5  <= '0';
            x6  <= '1';
            x7  <= '0';
            x8  <= '0';
            x9  <= '0';  
            
        when "01100100" => --t4q6
            x0  <= '0';
            x1  <= '0';
            x2  <= '1';
            x3  <= '0';
            x5  <= '0';
            x6  <= '1';
            x7  <= '0';
            x8  <= '0';
            x9  <= '0';   

        when "01100101" => --t5q6
            x0  <= '0';
            x1  <= '0';
            x2  <= '0';
            x3  <= '0';
            x5  <= '0';
            x6  <= '0';
            x7  <= '0';
            x8  <= '0';
            x9  <= '0'; 
            
        when "01100110" => --t6q6
            x0  <= '0';
            x1  <= '0';
            x2  <= '0';
            x3  <= '0';
            x5  <= '0';
            x6  <= '0';
            x7  <= '0';
            x8  <= '1';
            x9  <= '0'; 

        when "01100111" => --t7q6
            x0  <= '0';
            x1  <= '0';
            x2  <= '1';
            x3  <= '0';
            x5  <= '0';
            x6  <= '1';
            x7  <= '0';
            x8  <= '0';
            x9  <= '0'; 

        when "01101000" => --t8q6
            x0  <= '0';
            x1  <= '0';
            x2  <= '0';
            x3  <= '0';
            x5  <= '0';
            x6  <= '0';
            x7  <= '1';
            x8  <= '0';
            x9  <= '0'; 

        when "01101001" => --t9q6
            x0  <= '0';
            x1  <= '0';
            x2  <= '1';
            x3  <= '0';
            x5  <= '0';
            x6  <= '0';
            x7  <= '0';
            x8  <= '0';
            x9  <= '0'; 

        when "01101010" => --tAq6
            x0  <= '0';
            x1  <= '0';
            x2  <= '0';
            x3  <= '0';
            x5  <= '0';
            x6  <= '0';
            x7  <= '0';
            x8  <= '0';
            x9  <= '0'; 

        when "01101011" => --tBq6
            x0  <= '0';
            x1  <= '0';
            x2  <= '0';
            x3  <= '0';
            x5  <= '0';
            x6  <= '0';
            x7  <= '0';
            x8  <= '0';
            x9  <= '0'; 
------------  FIN -> 06h  AND A, [DIR]  

------------ 07h  OR A, [DIR]   
        --       q & t
        when "01110000" => --t0
            x0  <= '0';
            x1  <= '0';
            x2  <= '0';
            x3  <= '0';
            x5  <= '0';
            x6  <= '0';
            x7  <= '0';
            x8  <= '1';
            x9  <= '0';

        when "01110001" => --t1
            x0  <= '0';
            x1  <= '0';
            x2  <= '1';
            x3  <= '0';
            x5  <= '0';
            x6  <= '1';
            x7  <= '0';
            x8  <= '0';
            x9  <= '0';    
            
        when "01110010" => --t2
            x0  <= '1';
            x1  <= '0';
            x2  <= '0';
            x3  <= '0';
            x5  <= '0';
            x6  <= '0';
            x7  <= '0';
            x8  <= '0';
            x9  <= '0';    
            
        when "01110011" => --t3q7
            x0  <= '0';
            x1  <= '0';
            x2  <= '0';
            x3  <= '0';
            x5  <= '0';
            x6  <= '0';
            x7  <= '0';
            x8  <= '1';
            x9  <= '0';  
            
        when "01110100" => --t4q7
            x0  <= '0';
            x1  <= '0';
            x2  <= '1';
            x3  <= '0';
            x5  <= '0';
            x6  <= '1';
            x7  <= '0';
            x8  <= '0';
            x9  <= '0';   

        when "01110101" => --t5q7
            x0  <= '0';
            x1  <= '0';
            x2  <= '0';
            x3  <= '0';
            x5  <= '0';
            x6  <= '0';
            x7  <= '0';
            x8  <= '0';
            x9  <= '0'; 
            
        when "01110110" => --t6q7
            x0  <= '0';
            x1  <= '0';
            x2  <= '0';
            x3  <= '0';
            x5  <= '0';
            x6  <= '0';
            x7  <= '0';
            x8  <= '1';
            x9  <= '0'; 

        when "01110111" => --t7q7
            x0  <= '0';
            x1  <= '0';
            x2  <= '1';
            x3  <= '0';
            x5  <= '0';
            x6  <= '1';
            x7  <= '0';
            x8  <= '0';
            x9  <= '0'; 

        when "01111000" => --t8q7
            x0  <= '0';
            x1  <= '0';
            x2  <= '0';
            x3  <= '0';
            x5  <= '0';
            x6  <= '0';
            x7  <= '1';
            x8  <= '0';
            x9  <= '0'; 

        when "01111001" => --t9q7
            x0  <= '0';
            x1  <= '0';
            x2  <= '1';
            x3  <= '0';
            x5  <= '0';
            x6  <= '0';
            x7  <= '0';
            x8  <= '0';
            x9  <= '0'; 

        when "01111010" => --tAq7
            x0  <= '0';
            x1  <= '0';
            x2  <= '0';
            x3  <= '0';
            x5  <= '0';
            x6  <= '0';
            x7  <= '0';
            x8  <= '0';
            x9  <= '0'; 

        when "01111011" => --tBq7
            x0  <= '0';
            x1  <= '0';
            x2  <= '0';
            x3  <= '0';
            x5  <= '0';
            x6  <= '0';
            x7  <= '0';
            x8  <= '0';
            x9  <= '0'; 
------------  FIN -> 07h  OR A, [DIR]  

------------ 08h  JMP DIR   
        --       q & t
        when "10000000" => --t0
            x0  <= '0';
            x1  <= '0';
            x2  <= '0';
            x3  <= '0';
            x5  <= '0';
            x6  <= '0';
            x7  <= '0';
            x8  <= '1';
            x9  <= '0';

        when "10000001" => --t1
            x0  <= '0';
            x1  <= '0';
            x2  <= '1';
            x3  <= '0';
            x5  <= '0';
            x6  <= '1';
            x7  <= '0';
            x8  <= '0';
            x9  <= '0';    
            
        when "10000010" => --t2
            x0  <= '1';
            x1  <= '0';
            x2  <= '0';
            x3  <= '0';
            x5  <= '0';
            x6  <= '0';
            x7  <= '0';
            x8  <= '0';
            x9  <= '0';    
            
        when "10000011" => --t3q8
            x0  <= '0';
            x1  <= '0';
            x2  <= '0';
            x3  <= '0';
            x5  <= '0';
            x6  <= '0';
            x7  <= '0';
            x8  <= '1';
            x9  <= '0';  
            
        when "10000100" => --t4q8
            x0  <= '0';
            x1  <= '0';
            x2  <= '1';
            x3  <= '0';
            x5  <= '0';
            x6  <= '1';
            x7  <= '0';
            x8  <= '0';
            x9  <= '0';   

        when "10000101" => --t5q8
            x0  <= '0';
            x1  <= '0';
            x2  <= '0';
            x3  <= '0';
            x5  <= '0';
            x6  <= '0';
            x7  <= '0';
            x8  <= '0';
            x9  <= '0'; 
            
        when "10000110" => --t6q8
            x0  <= '0';
            x1  <= '0';
            x2  <= '0';
            x3  <= '0';
            x5  <= '0';
            x6  <= '0';
            x7  <= '0';
            x8  <= '1';
            x9  <= '0'; 

        when "10000111" => --t7q8
            x0  <= '0';
            x1  <= '0';
            x2  <= '1';
            x3  <= '0';
            x5  <= '0';
            x6  <= '1';
            x7  <= '0';
            x8  <= '0';
            x9  <= '0'; 

        when "10001000" => --t8q8
            x0  <= '0';
            x1  <= '0';
            x2  <= '0';
            x3  <= '0';
            x5  <= '1';
            x6  <= '0';
            x7  <= '0';
            x8  <= '0';
            x9  <= '0'; 

        when "10001001" => --t9q8
            x0  <= '0';
            x1  <= '0';
            x2  <= '0';
            x3  <= '0';
            x5  <= '0';
            x6  <= '0';
            x7  <= '0';
            x8  <= '0';
            x9  <= '0'; 

------------  FIN -> 08h  JMP [DIR]  

------------ 09h  JC DIR   
        --       q & t
        when "10010000" => --t0
            x0  <= '0';
            x1  <= '0';
            x2  <= '0';
            x3  <= '0';
            x5  <= '0';
            x6  <= '0';
            x7  <= '0';
            x8  <= '1';
            x9  <= '0';

        when "10010001" => --t1
            x0  <= '0';
            x1  <= '0';
            x2  <= '1';
            x3  <= '0';
            x5  <= '0';
            x6  <= '1';
            x7  <= '0';
            x8  <= '0';
            x9  <= '0';    
            
        when "10010010" => --t2
            x0  <= '1';
            x1  <= '0';
            x2  <= '0';
            x3  <= '0';
            x5  <= '0';
            x6  <= '0';
            x7  <= '0';
            x8  <= '0';
            x9  <= '0';    
            
        when "10010011" => --t3q9
            x0  <= '0';
            x1  <= '0';
            x2  <= '0';
            x3  <= '0';
            x5  <= '0';
            x6  <= '0';
            x7  <= '0';
            x8  <= '1';
            x9  <= '0';  
            
        when "10010100" => --t4q9
            x0  <= '0';
            x1  <= '0';
            x2  <= '1';
            x3  <= '0';
            x5  <= '0';
            x6  <= '1';
            x7  <= '0';
            x8  <= '0';
            x9  <= '0';   

        when "10010101" => --t5q9
            x0  <= '0';
            x1  <= '0';
            x2  <= '0';
            x3  <= '0';
            x5  <= '0';
            x6  <= '0';
            x7  <= '0';
            x8  <= '0';
            x9  <= '0'; 
            
        when "10010110" => --t6q9
            x0  <= '0';
            x1  <= '0';
            x2  <= '0';
            x3  <= '0';
            x5  <= '0';
            x6  <= '0';
            x7  <= '0';
            x8  <= '1';
            x9  <= '0'; 

        when "10010111" => --t7q9
            x0  <= '0';
            x1  <= '0';
            x2  <= '1';
            x3  <= '0';
            x5  <= '0';
            x6  <= '1';
            x7  <= '0';
            x8  <= '0';
            x9  <= '0'; 

        when "10011000" => --t8q9
           if (c_in = '1') then
                x0  <= '0';
                x1  <= '0';
                x2  <= '0';
                x3  <= '0';

                x5  <= '1';
                x6  <= '0';
                x7  <= '0';
                x8  <= '0';
                x9  <= '0';
 
            else
                x0  <= '0';
                x1  <= '0';
                x2  <= '0';
                x3  <= '0';

                x5  <= '0';
                x6  <= '0';
                x7  <= '0';
                x8  <= '0';
                x9  <= '0';

           end if ;

        when "10011001" => --t9q9
            x0  <= '0';
            x1  <= '0';
            x2  <= '0';
            x3  <= '0';
            x5  <= '0';
            x6  <= '0';
            x7  <= '0';
            x8  <= '0';
            x9  <= '0'; 

  
------------  FIN -> 09h  JC DIR    

------------ 0Ah  JZ DIR   
        --       q & t
        when "10100000" => --t0
            x0  <= '0';
            x1  <= '0';
            x2  <= '0';
            x3  <= '0';
            x5  <= '0';
            x6  <= '0';
            x7  <= '0';
            x8  <= '1';
            x9  <= '0';

        when "10100001" => --t1
            x0  <= '0';
            x1  <= '0';
            x2  <= '1';
            x3  <= '0';
            x5  <= '0';
            x6  <= '1';
            x7  <= '0';
            x8  <= '0';
            x9  <= '0';    
            
        when "10100010" => --t2
            x0  <= '1';
            x1  <= '0';
            x2  <= '0';
            x3  <= '0';
            x5  <= '0';
            x6  <= '0';
            x7  <= '0';
            x8  <= '0';
            x9  <= '0';    
            
        when "10100011" => --t3qA
            x0  <= '0';
            x1  <= '0';
            x2  <= '0';
            x3  <= '0';
            x5  <= '0';
            x6  <= '0';
            x7  <= '0';
            x8  <= '1';
            x9  <= '0';  
            
        when "10100100" => --t4qA
            x0  <= '0';
            x1  <= '0';
            x2  <= '1';
            x3  <= '0';
            x5  <= '0';
            x6  <= '1';
            x7  <= '0';
            x8  <= '0';
            x9  <= '0';   

        when "10100101" => --t5qA
            x0  <= '0';
            x1  <= '0';
            x2  <= '0';
            x3  <= '0';
            x5  <= '0';
            x6  <= '0';
            x7  <= '0';
            x8  <= '0';
            x9  <= '0'; 
            
        when "10100110" => --t6qA
            x0  <= '0';
            x1  <= '0';
            x2  <= '0';
            x3  <= '0';
            x5  <= '0';
            x6  <= '0';
            x7  <= '0';
            x8  <= '1';
            x9  <= '0'; 

        when "10100111" => --t7qA
            x0  <= '0';
            x1  <= '0';
            x2  <= '1';
            x3  <= '0';
            x5  <= '0';
            x6  <= '1';
            x7  <= '0';
            x8  <= '0';
            x9  <= '0'; 

        when "10101000" => --t8qA
           if (z_in = '1') then
                x0  <= '0';
                x1  <= '0';
                x2  <= '0';
                x3  <= '0';

                x5  <= '1';
                x6  <= '0';
                x7  <= '0';
                x8  <= '0';
                x9  <= '0';
 
            else
                x0  <= '0';
                x1  <= '0';
                x2  <= '0';
                x3  <= '0';

                x5  <= '0';
                x6  <= '0';
                x7  <= '0';
                x8  <= '0';
                x9  <= '0';
 
           end if ;

        when "10101001" => --t9qA
            x0  <= '0';
            x1  <= '0';
            x2  <= '0';
            x3  <= '0';
            x5  <= '0';
            x6  <= '0';
            x7  <= '0';
            x8  <= '0';
            x9  <= '0'; 

  
------------  FIN -> 0Ah  JZ DIR  

------------ 0Bh  JSR DIR   
        --       q & t
        when "10110000" => --t0
            x0  <= '0';
            x1  <= '0';
            x2  <= '0';
            x3  <= '0';
            x5  <= '0';
            x6  <= '0';
            x7  <= '0';
            x8  <= '1';
            x9  <= '0';

        when "10110001" => --t1
            x0  <= '0';
            x1  <= '0';
            x2  <= '1';
            x3  <= '0';
            x5  <= '0';
            x6  <= '1';
            x7  <= '0';
            x8  <= '0';
            x9  <= '0';    
            
        when "10110010" => --t2
            x0  <= '1';
            x1  <= '0';
            x2  <= '0';
            x3  <= '0';
            x5  <= '0';
            x6  <= '0';
            x7  <= '0';
            x8  <= '0';
            x9  <= '0';    
            
        when "10110011" => --t3qB
            x0  <= '0';
            x1  <= '0';
            x2  <= '0';
            x3  <= '0';
            x5  <= '0';
            x6  <= '0';
            x7  <= '0';
            x8  <= '1';
            x9  <= '0';  
            
        when "10110100" => --t4qB
            x0  <= '0';
            x1  <= '0';
            x2  <= '1';
            x3  <= '0';
            x5  <= '0';
            x6  <= '1';
            x7  <= '0';
            x8  <= '0';
            x9  <= '0';   

        when "10110101" => --t5qB
            x0  <= '0';
            x1  <= '0';
            x2  <= '0';
            x3  <= '0';
            x5  <= '0';
            x6  <= '0';
            x7  <= '0';
            x8  <= '1';
            x9  <= '0'; 
            
        when "10110110" => --t6qB
            x0  <= '0';
            x1  <= '0';
            x2  <= '1';
            x3  <= '0';
            x5  <= '0';
            x6  <= '1';
            x7  <= '0';
            x8  <= '0';
            x9  <= '0'; 

        when "10110111" => --t7qB
            x0  <= '0';
            x1  <= '0';
            x2  <= '0';
            x3  <= '0';
            x5  <= '0';
            x6  <= '0';
            x7  <= '0';
            x8  <= '0';
            x9  <= '1'; 

        when "10111000" => --t8qB
                x0  <= '0';
                x1  <= '0';
                x2  <= '0';
                x3  <= '1';

                x5  <= '0';
                x6  <= '0';
                x7  <= '0';
                x8  <= '0';
                x9  <= '0';

        when "10111001" => --t9qB
            x0  <= '0';
            x1  <= '0';
            x2  <= '0';
            x3  <= '0';
            x5  <= '0';
            x6  <= '0';
            x7  <= '0';
            x8  <= '0';
            x9  <= '0'; 

        when "10111010" => --tAqB
            x0  <= '0';
            x1  <= '0';
            x2  <= '0';
            x3  <= '0';
            x5  <= '0';
            x6  <= '0';
            x7  <= '0';
            x8  <= '0';
            x9  <= '1'; 
  
        when "10111011" => --tBqB
            x0  <= '0';
            x1  <= '0';
            x2  <= '0';
            x3  <= '0';
            x5  <= '0';
            x6  <= '0';
            x7  <= '0';
            x8  <= '0';
            x9  <= '0';
            
        when "10111100" => --tCqB
            x0  <= '0';
            x1  <= '0';
            x2  <= '0';
            x3  <= '0';
            x5  <= '0';
            x6  <= '0';
            x7  <= '0';
            x8  <= '0';
            x9  <= '0';
            
        when "10111101" => --tDqB
            x0  <= '0';
            x1  <= '1';
            x2  <= '0';
            x3  <= '0';
            x5  <= '0';
            x6  <= '0';
            x7  <= '0';
            x8  <= '0';
            x9  <= '0'; 

        when "10111110" => --tEqB
            x0  <= '0';
            x1  <= '0';
            x2  <= '0';
            x3  <= '0';
            x5  <= '1';
            x6  <= '0';
            x7  <= '0';
            x8  <= '0';
            x9  <= '0'; 

        when "10111111" => --tFqB
            x0  <= '0';
            x1  <= '0';
            x2  <= '0';
            x3  <= '0';
            x5  <= '0';
            x6  <= '0';
            x7  <= '0';
            x8  <= '0';
            x9  <= '0'; 
------------  FIN -> 0Bh  JSR DIR  

------------ 0Ch  RTS 
        --       q & t
        when "11000000" => --t0
            x0  <= '0';
            x1  <= '0';
            x2  <= '0';
            x3  <= '0';
            x5  <= '0';
            x6  <= '0';
            x7  <= '0';
            x8  <= '1';
            x9  <= '0';

        when "11000001" => --t1
            x0  <= '0';
            x1  <= '0';
            x2  <= '1';
            x3  <= '0';
            x5  <= '0';
            x6  <= '1';
            x7  <= '0';
            x8  <= '0';
            x9  <= '0';    
            
        when "11000010" => --t2
            x0  <= '1';
            x1  <= '0';
            x2  <= '0';
            x3  <= '0';
            x5  <= '0';
            x6  <= '0';
            x7  <= '0';
            x8  <= '0';
            x9  <= '0';    
            
        when "11000011" => --t3qC
            x0  <= '0';
            x1  <= '0';
            x2  <= '0';
            x3  <= '0';
            x5  <= '0';
            x6  <= '0';
            x7  <= '0';
            x8  <= '0';
            x9  <= '0';  
            
        when "11000100" => --t4qC
            x0  <= '0';
            x1  <= '0';
            x2  <= '0';
            x3  <= '0';
            x5  <= '0';
            x6  <= '0';
            x7  <= '0';
            x8  <= '0';
            x9  <= '1';   

        when "11000101" => --t5qC
            x0  <= '0';
            x1  <= '0';
            x2  <= '1';
            x3  <= '0';
            x5  <= '0';
            x6  <= '0';
            x7  <= '0';
            x8  <= '1';
            x9  <= '0'; 
            
        when "11000110" => --t6qC
            x0  <= '0';
            x1  <= '0';
            x2  <= '0';
            x3  <= '0';
            x5  <= '0';
            x6  <= '0';
            x7  <= '0';
            x8  <= '0';
            x9  <= '0'; 

        when "11000111" => --t7qC
            x0  <= '0';
            x1  <= '0';
            x2  <= '0';
            x3  <= '0';
            x5  <= '0';
            x6  <= '0';
            x7  <= '0';
            x8  <= '0';
            x9  <= '1'; 

        when "11001000" => --t8qC
                x0  <= '0';
                x1  <= '0';
                x2  <= '1';
                x3  <= '0';
                x5  <= '0';
                x6  <= '0';
                x7  <= '0';
                x8  <= '0';
                x9  <= '1';

        when "11001001" => --t9qC
            x0  <= '0';
            x1  <= '0';
            x2  <= '0';
            x3  <= '0';
            x5  <= '1';
            x6  <= '0';
            x7  <= '0';
            x8  <= '0';
            x9  <= '0'; 

        when "11001010" => --tAqC
            x0  <= '0';
            x1  <= '0';
            x2  <= '0';
            x3  <= '0';
            x5  <= '0';
            x6  <= '0';
            x7  <= '0';
            x8  <= '0';
            x9  <= '0'; 
------------  FIN -> 0Ch  RTS  

------------  0Dh  LSL A 
        --       q & t
        when "11010000" => --t0
            x0  <= '0';
            x1  <= '0';
            x2  <= '0';
            x3  <= '0';
            x5  <= '0';
            x6  <= '0';
            x7  <= '0';
            x8  <= '1';
            x9  <= '0';

        when "11010001" => --t1
            x0  <= '0';
            x1  <= '0';
            x2  <= '1';
            x3  <= '0';
            x5  <= '0';
            x6  <= '1';
            x7  <= '0';
            x8  <= '0';
            x9  <= '0';    
            
        when "11010010" => --t2
            x0  <= '1';
            x1  <= '0';
            x2  <= '0';
            x3  <= '0';
            x5  <= '0';
            x6  <= '0';
            x7  <= '0';
            x8  <= '0';
            x9  <= '0';    
            
        when "11010011" => --t3qD
            x0  <= '0';
            x1  <= '0';
            x2  <= '0';
            x3  <= '0';
            x5  <= '0';
            x6  <= '0';
            x7  <= '0';
            x8  <= '0';
            x9  <= '0';  
            
        when "11010100" => --t4qD
            x0  <= '0';
            x1  <= '0';
            x2  <= '0';
            x3  <= '0';
            x5  <= '0';
            x6  <= '0';
            x7  <= '0';
            x8  <= '0';
            x9  <= '0';   
------------  FIN -> 0Dh  LSL A  


------------  0Eh  LSR A 
        --       q & t
        when "11100000" => --t0
            x0  <= '0';
            x1  <= '0';
            x2  <= '0';
            x3  <= '0';
            x5  <= '0';
            x6  <= '0';
            x7  <= '0';
            x8  <= '1';
            x9  <= '0';

        when "11100001" => --t1
            x0  <= '0';
            x1  <= '0';
            x2  <= '1';
            x3  <= '0';
            x5  <= '0';
            x6  <= '1';
            x7  <= '0';
            x8  <= '0';
            x9  <= '0';    
            
        when "11100010" => --t2
            x0  <= '1';
            x1  <= '0';
            x2  <= '0';
            x3  <= '0';
            x5  <= '0';
            x6  <= '0';
            x7  <= '0';
            x8  <= '0';
            x9  <= '0';    
            
        when "11100011" => --t3qE
            x0  <= '0';
            x1  <= '0';
            x2  <= '0';
            x3  <= '0';
            x5  <= '0';
            x6  <= '0';
            x7  <= '0';
            x8  <= '0';
            x9  <= '0';  
            
        when "11100100" => --t4qE
            x0  <= '0';
            x1  <= '0';
            x2  <= '0';
            x3  <= '0';
            x5  <= '0';
            x6  <= '0';
            x7  <= '0';
            x8  <= '0';
            x9  <= '0';   
------------  FIN -> 0Eh  LSR A  

------------  0Eh  NOT A 
        --       q & t
        when "11110000" => --t0
            x0  <= '0';
            x1  <= '0';
            x2  <= '0';
            x3  <= '0';
            x5  <= '0';
            x6  <= '0';
            x7  <= '0';
            x8  <= '1';
            x9  <= '0';

        when "11110001" => --t1
            x0  <= '0';
            x1  <= '0';
            x2  <= '1';
            x3  <= '0';
            x5  <= '0';
            x6  <= '1';
            x7  <= '0';
            x8  <= '0';
            x9  <= '0';    
            
        when "11110010" => --t2
            x0  <= '1';
            x1  <= '0';
            x2  <= '0';
            x3  <= '0';
            x5  <= '0';
            x6  <= '0';
            x7  <= '0';
            x8  <= '0';
            x9  <= '0';    
            
        when "11110011" => --t3qF
            x0  <= '0';
            x1  <= '0';
            x2  <= '0';
            x3  <= '0';
            x5  <= '0';
            x6  <= '0';
            x7  <= '0';
            x8  <= '0';
            x9  <= '0';  
            
        when "11110100" => --t4qF
            x0  <= '0';
            x1  <= '0';
            x2  <= '0';
            x3  <= '0';
            x5  <= '0';
            x6  <= '0';
            x7  <= '0';
            x8  <= '0';
            x9  <= '0';   
------------  FIN -> 0Fh  NOT A  
when others => -- reset
            x0  <= '0';
            x1  <= '0';
            x2  <= '0';
            x3  <= '0';
            x5  <= '0';
            x6  <= '0';
            x7  <= '0';
            x8  <= '0';
            x9  <= '0';   
        end case ;
           
    end process;
   Xs_out <= x9 & x8 & x7 & x6 & x5 & x3 & x2 & x1 & & x0 ;
end architecture ;


