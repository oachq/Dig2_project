library ieee ;
    use ieee.std_logic_1164.all ;
    use ieee.numeric_std.all ;
    use IEEE.std_logic_arith.all;
    use IEEE.std_logic_unsigned.all;

entity UC is
    generic (
        wl_Q:   integer:= 4;
        wl_T:   integer:= 4;
        wl_Xs:  integer:= 20
    );
  port (
    q_in:   in  std_logic_vector(wl_Q-1 downto 0);
    t_in:   in  std_logic_vector(wl_T-1 downto 0);
    c_in:   in  std_logic;
    z_in:   in  std_logic;
    Xs_out: out std_logic_vector(wl_Xs downto 0)
  ) ;
end UC ; 
--:= (others => '0' )
architecture arch of UC is

    signal control : std_logic_vector(8 downto 0);  -- control de entradas
    signal xs: std_logic_vector(wl_Xs downto 0); -- array salida xs
    signal flags: std_logic_vector(1 downto 0);-- entradas banderas
begin
    
   control <= q_in & t_in; -- concatenando entradas q y t

    process (q_in, t_in, control )
    begin
        case( control ) is
------------  00h  MOV A, N
        --       q & t
            when "0000"&"0000" => --t0
                xs(0)  <= '0';
                xs(1)  <= '0';
                xs(2)  <= '0';
                xs(3)  <= '0';
                xs(4)  <= '0';
                xs(5)  <= '0';
                xs(6)  <= '0';
                xs(7)  <= '0';
                xs(8)  <= '1';
                xs(9)  <= '0';
                xs(10) <= '0';
                xs(11) <= '0';
                xs(12) <= '0';
                xs(13) <= '0';
                xs(14) <= '0';
                xs(15) <= '0';
                xs(16) <= '0';
                xs(17) <= '0';
                xs(18) <= '0';
                xs(19) <= '0';
                xs(20) <= '0';

            when "0000"&"0001" => --t1
                xs(0)  <= '0';
                xs(1)  <= '0';
                xs(2)  <= '1';
                xs(3)  <= '0';
                xs(4)  <= '0';
                xs(5)  <= '0';
                xs(6)  <= '1';
                xs(7)  <= '0';
                xs(8)  <= '0';
                xs(9)  <= '0';
                xs(10) <= '0';
                xs(11) <= '0';
                xs(12) <= '0';
                xs(13) <= '0';
                xs(14) <= '0';
                xs(15) <= '0';
                xs(16) <= '0';
                xs(17) <= '0';
                xs(18) <= '0';
                xs(19) <= '0';
                xs(20) <= '0';    
                
            when "0000"&"0010" => --t2
                xs(0)  <= '1';
                xs(1)  <= '0';
                xs(2)  <= '0';
                xs(3)  <= '0';
                xs(4)  <= '0';
                xs(5)  <= '0';
                xs(6)  <= '0';
                xs(7)  <= '0';
                xs(8)  <= '0';
                xs(9)  <= '0';
                xs(10) <= '0';
                xs(11) <= '0';
                xs(12) <= '0';
                xs(13) <= '0';
                xs(14) <= '0';
                xs(15) <= '0';
                xs(16) <= '0';
                xs(17) <= '0';
                xs(18) <= '0';
                xs(19) <= '0';
                xs(20) <= '0';    
                
            when "0000"&"0011" => --t3q0
                xs(0)  <= '0';
                xs(1)  <= '0';
                xs(2)  <= '0';
                xs(3)  <= '0';
                xs(4)  <= '0';
                xs(5)  <= '0';
                xs(6)  <= '0';
                xs(7)  <= '0';
                xs(8)  <= '1';
                xs(9)  <= '0';
                xs(10) <= '0';
                xs(11) <= '0';
                xs(12) <= '0';
                xs(13) <= '0';
                xs(14) <= '0';
                xs(15) <= '0';
                xs(16) <= '0';
                xs(17) <= '0';
                xs(18) <= '0';
                xs(19) <= '0';
                xs(20) <= '0';  
                
            when "0000"&"0100" => --t4q0
                xs(0)  <= '0';
                xs(1)  <= '0';
                xs(2)  <= '1';
                xs(3)  <= '0';
                xs(4)  <= '0';
                xs(5)  <= '0';
                xs(6)  <= '1';
                xs(7)  <= '0';
                xs(8)  <= '0';
                xs(9)  <= '0';
                xs(10) <= '0';
                xs(11) <= '0';
                xs(12) <= '0';
                xs(13) <= '0';
                xs(14) <= '0';
                xs(15) <= '0';
                xs(16) <= '0';
                xs(17) <= '0';
                xs(18) <= '0';
                xs(19) <= '0';
                xs(20) <= '0';   

            when "0000"&"0101" => --t5q0
                xs(0)  <= '0';
                xs(1)  <= '0';
                xs(2)  <= '0';
                xs(3)  <= '0';
                xs(4)  <= '0';
                xs(5)  <= '0';
                xs(6)  <= '0';
                xs(7)  <= '0';
                xs(8)  <= '0';
                xs(9)  <= '0';
                xs(10) <= '0';
                xs(11) <= '0';
                xs(12) <= '0';
                xs(13) <= '0';
                xs(14) <= '0';
                xs(15) <= '1';
                xs(16) <= '1';
                xs(17) <= '1';
                xs(18) <= '0';
                xs(19) <= '1';
                xs(20) <= '0'; 
            
            when "0000"&"0110" => --t6q0
                xs(0)  <= '0';
                xs(1)  <= '0';
                xs(2)  <= '0';
                xs(3)  <= '0';
                xs(4)  <= '0';
                xs(5)  <= '0';
                xs(6)  <= '0';
                xs(7)  <= '0';
                xs(8)  <= '0';
                xs(9)  <= '0';
                xs(10) <= '0';
                xs(11) <= '0';
                xs(12) <= '0';
                xs(13) <= '0';
                xs(14) <= '1';
                xs(15) <= '0';
                xs(16) <= '0';
                xs(17) <= '0';
                xs(18) <= '0';
                xs(19) <= '0';
                xs(20) <= '0';         
------------  FIN -> 00h  MOV A, N            
            
------------  01h  MOV A, [DIR]
        --       q & t
            when "0001"&"0000" => --t0
                xs(0)  <= '0';
                xs(1)  <= '0';
                xs(2)  <= '0';
                xs(3)  <= '0';
                xs(4)  <= '0';
                xs(5)  <= '0';
                xs(6)  <= '0';
                xs(7)  <= '0';
                xs(8)  <= '1';
                xs(9)  <= '0';
                xs(10) <= '0';
                xs(11) <= '0';
                xs(12) <= '0';
                xs(13) <= '0';
                xs(14) <= '0';
                xs(15) <= '0';
                xs(16) <= '0';
                xs(17) <= '0';
                xs(18) <= '0';
                xs(19) <= '0';
                xs(20) <= '0';

            when "0001"&"0001" => --t1
                xs(0)  <= '0';
                xs(1)  <= '0';
                xs(2)  <= '1';
                xs(3)  <= '0';
                xs(4)  <= '0';
                xs(5)  <= '0';
                xs(6)  <= '1';
                xs(7)  <= '0';
                xs(8)  <= '0';
                xs(9)  <= '0';
                xs(10) <= '0';
                xs(11) <= '0';
                xs(12) <= '0';
                xs(13) <= '0';
                xs(14) <= '0';
                xs(15) <= '0';
                xs(16) <= '0';
                xs(17) <= '0';
                xs(18) <= '0';
                xs(19) <= '0';
                xs(20) <= '0';    

            when "0001"&"0010" => --t2
                xs(0)  <= '1';
                xs(1)  <= '0';
                xs(2)  <= '0';
                xs(3)  <= '0';
                xs(4)  <= '0';
                xs(5)  <= '0';
                xs(6)  <= '0';
                xs(7)  <= '0';
                xs(8)  <= '0';
                xs(9)  <= '0';
                xs(10) <= '0';
                xs(11) <= '0';
                xs(12) <= '0';
                xs(13) <= '0';
                xs(14) <= '0';
                xs(15) <= '0';
                xs(16) <= '0';
                xs(17) <= '0';
                xs(18) <= '0';
                xs(19) <= '0';
                xs(20) <= '0';    

            when "0001"&"0011" => --t3q1
                xs(0)  <= '0';
                xs(1)  <= '0';
                xs(2)  <= '0';
                xs(3)  <= '0';
                xs(4)  <= '0';
                xs(5)  <= '0';
                xs(6)  <= '0';
                xs(7)  <= '0';
                xs(8)  <= '1';
                xs(9)  <= '0';
                xs(10) <= '0';
                xs(11) <= '0';
                xs(12) <= '0';
                xs(13) <= '0';
                xs(14) <= '0';
                xs(15) <= '0';
                xs(16) <= '0';
                xs(17) <= '0';
                xs(18) <= '0';
                xs(19) <= '0';
                xs(20) <= '0';  

            when "0001"&"0100" => --t4q1
                xs(0)  <= '0';
                xs(1)  <= '0';
                xs(2)  <= '1';
                xs(3)  <= '0';
                xs(4)  <= '0';
                xs(5)  <= '0';
                xs(6)  <= '1';
                xs(7)  <= '0';
                xs(8)  <= '0';
                xs(9)  <= '0';
                xs(10) <= '0';
                xs(11) <= '0';
                xs(12) <= '0';
                xs(13) <= '0';
                xs(14) <= '0';
                xs(15) <= '0';
                xs(16) <= '0';
                xs(17) <= '0';
                xs(18) <= '0';
                xs(19) <= '0';
                xs(20) <= '0';   

            when "0001"&"0101" => --t5q1
                xs(0)  <= '0';
                xs(1)  <= '0';
                xs(2)  <= '0';
                xs(3)  <= '0';
                xs(4)  <= '0';
                xs(5)  <= '0';
                xs(6)  <= '0';
                xs(7)  <= '0';
                xs(8)  <= '0';
                xs(9)  <= '0';
                xs(10) <= '1';
                xs(11) <= '0';
                xs(12) <= '0';
                xs(13) <= '0';
                xs(14) <= '0';
                xs(15) <= '0';
                xs(16) <= '0';
                xs(17) <= '0';
                xs(18) <= '0';
                xs(19) <= '0';
                xs(20) <= '0'; 

            when "0001"&"0110" => --t6q1
                xs(0)  <= '0';
                xs(1)  <= '0';
                xs(2)  <= '0';
                xs(3)  <= '0';
                xs(4)  <= '0';
                xs(5)  <= '0';
                xs(6)  <= '0';
                xs(7)  <= '0';
                xs(8)  <= '1';
                xs(9)  <= '0';
                xs(10) <= '0';
                xs(11) <= '0';
                xs(12) <= '0';
                xs(13) <= '0';
                xs(14) <= '0';
                xs(15) <= '0';
                xs(16) <= '0';
                xs(17) <= '0';
                xs(18) <= '0';
                xs(19) <= '0';
                xs(20) <= '0';
                
            when "0001"&"0111" => --t7q1
                xs(0)  <= '0';
                xs(1)  <= '0';
                xs(2)  <= '1';
                xs(3)  <= '0';
                xs(4)  <= '0';
                xs(5)  <= '0';
                xs(6)  <= '1';
                xs(7)  <= '0';
                xs(8)  <= '0';
                xs(9)  <= '0';
                xs(10) <= '0';
                xs(11) <= '0';
                xs(12) <= '0';
                xs(13) <= '0';
                xs(14) <= '0';
                xs(15) <= '0';
                xs(16) <= '0';
                xs(17) <= '0';
                xs(18) <= '0';
                xs(19) <= '0';
                xs(20) <= '0';
                
            when "0001"&"1000" => --t8q1
                xs(0)  <= '0';
                xs(1)  <= '0';
                xs(2)  <= '0';
                xs(3)  <= '0';
                xs(4)  <= '0';
                xs(5)  <= '0';
                xs(6)  <= '0';
                xs(7)  <= '1';
                xs(8)  <= '0';
                xs(9)  <= '0';
                xs(10) <= '0';
                xs(11) <= '0';
                xs(12) <= '0';
                xs(13) <= '0';
                xs(14) <= '0';
                xs(15) <= '0';
                xs(16) <= '0';
                xs(17) <= '0';
                xs(18) <= '0';
                xs(19) <= '0';
                xs(20) <= '0';
                
            when "0001"&"1001" => --t9q1
                xs(0)  <= '0';
                xs(1)  <= '0';
                xs(2)  <= '1';
                xs(3)  <= '0';
                xs(4)  <= '0';
                xs(5)  <= '0';
                xs(6)  <= '0';
                xs(7)  <= '0';
                xs(8)  <= '0';
                xs(9)  <= '0';
                xs(10) <= '0';
                xs(11) <= '0';
                xs(12) <= '0';
                xs(13) <= '0';
                xs(14) <= '0';
                xs(15) <= '0';
                xs(16) <= '0';
                xs(17) <= '0';
                xs(18) <= '0';
                xs(19) <= '0';
                xs(20) <= '0';  
                
            when "0001"&"1010" => --tAq1 
                xs(0)  <= '0';
                xs(1)  <= '0';
                xs(2)  <= '0';
                xs(3)  <= '0';
                xs(4)  <= '0';
                xs(5)  <= '0';
                xs(6)  <= '0';
                xs(7)  <= '0';
                xs(8)  <= '0';
                xs(9)  <= '0';
                xs(10) <= '0';
                xs(11) <= '0';
                xs(12) <= '0';
                xs(13) <= '0';
                xs(14) <= '0';
                xs(15) <= '1';
                xs(16) <= '1';
                xs(17) <= '1';
                xs(18) <= '0';
                xs(19) <= '1';
                xs(20) <= '0';

            when "0001"&"1011" => --tBq1
                xs(0)  <= '0';
                xs(1)  <= '0';
                xs(2)  <= '0';
                xs(3)  <= '0';
                xs(4)  <= '0';
                xs(5)  <= '0';
                xs(6)  <= '0';
                xs(7)  <= '0';
                xs(8)  <= '0';
                xs(9)  <= '0';
                xs(10) <= '0';
                xs(11) <= '0';
                xs(12) <= '0';
                xs(13) <= '0';
                xs(14) <= '1';
                xs(15) <= '0';
                xs(16) <= '0';
                xs(17) <= '0';
                xs(18) <= '0';
                xs(19) <= '0';
                xs(20) <= '0';
------------  FIN -> MOV A, [DIR]           
    
------------ 02h  MOV SP, [N]
        --       q & t
        when "0010"&"0000" => --t0
            xs(0)  <= '0';
            xs(1)  <= '0';
            xs(2)  <= '0';
            xs(3)  <= '0';
            xs(4)  <= '0';
            xs(5)  <= '0';
            xs(6)  <= '0';
            xs(7)  <= '0';
            xs(8)  <= '1';
            xs(9)  <= '0';
            xs(10) <= '0';
            xs(11) <= '0';
            xs(12) <= '0';
            xs(13) <= '0';
            xs(14) <= '0';
            xs(15) <= '0';
            xs(16) <= '0';
            xs(17) <= '0';
            xs(18) <= '0';
            xs(19) <= '0';
            xs(20) <= '0';

        when "0010"&"0001" => --t1
            xs(0)  <= '0';
            xs(1)  <= '0';
            xs(2)  <= '1';
            xs(3)  <= '0';
            xs(4)  <= '0';
            xs(5)  <= '0';
            xs(6)  <= '1';
            xs(7)  <= '0';
            xs(8)  <= '0';
            xs(9)  <= '0';
            xs(10) <= '0';
            xs(11) <= '0';
            xs(12) <= '0';
            xs(13) <= '0';
            xs(14) <= '0';
            xs(15) <= '0';
            xs(16) <= '0';
            xs(17) <= '0';
            xs(18) <= '0';
            xs(19) <= '0';
            xs(20) <= '0';    
            
        when "0010"&"0010" => --t2
            xs(0)  <= '1';
            xs(1)  <= '0';
            xs(2)  <= '0';
            xs(3)  <= '0';
            xs(4)  <= '0';
            xs(5)  <= '0';
            xs(6)  <= '0';
            xs(7)  <= '0';
            xs(8)  <= '0';
            xs(9)  <= '0';
            xs(10) <= '0';
            xs(11) <= '0';
            xs(12) <= '0';
            xs(13) <= '0';
            xs(14) <= '0';
            xs(15) <= '0';
            xs(16) <= '0';
            xs(17) <= '0';
            xs(18) <= '0';
            xs(19) <= '0';
            xs(20) <= '0';    
            
        when "0010"&"0011" => --t3q2
            xs(0)  <= '0';
            xs(1)  <= '0';
            xs(2)  <= '0';
            xs(3)  <= '0';
            xs(4)  <= '0';
            xs(5)  <= '0';
            xs(6)  <= '0';
            xs(7)  <= '0';
            xs(8)  <= '1';
            xs(9)  <= '0';
            xs(10) <= '0';
            xs(11) <= '0';
            xs(12) <= '0';
            xs(13) <= '0';
            xs(14) <= '0';
            xs(15) <= '0';
            xs(16) <= '0';
            xs(17) <= '0';
            xs(18) <= '0';
            xs(19) <= '0';
            xs(20) <= '0';  
            
        when "0010"&"0100" => --t4q2
            xs(0)  <= '0';
            xs(1)  <= '0';
            xs(2)  <= '1';
            xs(3)  <= '0';
            xs(4)  <= '0';
            xs(5)  <= '0';
            xs(6)  <= '1';
            xs(7)  <= '0';
            xs(8)  <= '0';
            xs(9)  <= '0';
            xs(10) <= '0';
            xs(11) <= '0';
            xs(12) <= '0';
            xs(13) <= '0';
            xs(14) <= '0';
            xs(15) <= '0';
            xs(16) <= '0';
            xs(17) <= '0';
            xs(18) <= '0';
            xs(19) <= '0';
            xs(20) <= '0';   

        when "0010"&"0101" => --t5q2
            xs(0)  <= '0';
            xs(1)  <= '0';
            xs(2)  <= '0';
            xs(3)  <= '0';
            xs(4)  <= '0';
            xs(5)  <= '0';
            xs(6)  <= '0';
            xs(7)  <= '0';
            xs(8)  <= '0';
            xs(9)  <= '0';
            xs(10) <= '0';
            xs(11) <= '1';
            xs(12) <= '0';
            xs(13) <= '0';
            xs(14) <= '0';
            xs(15) <= '0';
            xs(16) <= '0';
            xs(17) <= '0';
            xs(18) <= '0';
            xs(19) <= '0';
            xs(20) <= '0'; 
            
        when "0010"&"0110" => --t6q2
            xs(0)  <= '0';
            xs(1)  <= '0';
            xs(2)  <= '0';
            xs(3)  <= '0';
            xs(4)  <= '0';
            xs(5)  <= '0';
            xs(6)  <= '0';
            xs(7)  <= '0';
            xs(8)  <= '0';
            xs(9)  <= '0';
            xs(10) <= '0';
            xs(11) <= '0';
            xs(12) <= '0';
            xs(13) <= '0';
            xs(14) <= '1';
            xs(15) <= '0';
            xs(16) <= '0';
            xs(17) <= '0';
            xs(18) <= '0';
            xs(19) <= '0';
            xs(20) <= '0';         
------------  FIN -> 02h  MOV SP, [N]           
            
------------ 03h  MOV [DIR], A
        --       q & t
        when "0011"&"0000" => --t0
            xs(0)  <= '0';
            xs(1)  <= '0';
            xs(2)  <= '0';
            xs(3)  <= '0';
            xs(4)  <= '0';
            xs(5)  <= '0';
            xs(6)  <= '0';
            xs(7)  <= '0';
            xs(8)  <= '1';
            xs(9)  <= '0';
            xs(10) <= '0';
            xs(11) <= '0';
            xs(12) <= '0';
            xs(13) <= '0';
            xs(14) <= '0';
            xs(15) <= '0';
            xs(16) <= '0';
            xs(17) <= '0';
            xs(18) <= '0';
            xs(19) <= '0';
            xs(20) <= '0';

        when "0011"&"0001" => --t1
            xs(0)  <= '0';
            xs(1)  <= '0';
            xs(2)  <= '1';
            xs(3)  <= '0';
            xs(4)  <= '0';
            xs(5)  <= '0';
            xs(6)  <= '1';
            xs(7)  <= '0';
            xs(8)  <= '0';
            xs(9)  <= '0';
            xs(10) <= '0';
            xs(11) <= '0';
            xs(12) <= '0';
            xs(13) <= '0';
            xs(14) <= '0';
            xs(15) <= '0';
            xs(16) <= '0';
            xs(17) <= '0';
            xs(18) <= '0';
            xs(19) <= '0';
            xs(20) <= '0';    
            
        when "0011"&"0010" => --t2
            xs(0)  <= '1';
            xs(1)  <= '0';
            xs(2)  <= '0';
            xs(3)  <= '0';
            xs(4)  <= '0';
            xs(5)  <= '0';
            xs(6)  <= '0';
            xs(7)  <= '0';
            xs(8)  <= '0';
            xs(9)  <= '0';
            xs(10) <= '0';
            xs(11) <= '0';
            xs(12) <= '0';
            xs(13) <= '0';
            xs(14) <= '0';
            xs(15) <= '0';
            xs(16) <= '0';
            xs(17) <= '0';
            xs(18) <= '0';
            xs(19) <= '0';
            xs(20) <= '0';    
            
        when "0011"&"0011" => --t3q3
            xs(0)  <= '0';
            xs(1)  <= '0';
            xs(2)  <= '0';
            xs(3)  <= '0';
            xs(4)  <= '0';
            xs(5)  <= '0';
            xs(6)  <= '0';
            xs(7)  <= '0';
            xs(8)  <= '1';
            xs(9)  <= '0';
            xs(10) <= '0';
            xs(11) <= '0';
            xs(12) <= '0';
            xs(13) <= '0';
            xs(14) <= '0';
            xs(15) <= '0';
            xs(16) <= '0';
            xs(17) <= '0';
            xs(18) <= '0';
            xs(19) <= '0';
            xs(20) <= '0';  
            
        when "0011"&"0100" => --t4q3
            xs(0)  <= '0';
            xs(1)  <= '0';
            xs(2)  <= '1';
            xs(3)  <= '0';
            xs(4)  <= '0';
            xs(5)  <= '0';
            xs(6)  <= '1';
            xs(7)  <= '0';
            xs(8)  <= '0';
            xs(9)  <= '0';
            xs(10) <= '0';
            xs(11) <= '0';
            xs(12) <= '0';
            xs(13) <= '0';
            xs(14) <= '0';
            xs(15) <= '0';
            xs(16) <= '0';
            xs(17) <= '0';
            xs(18) <= '0';
            xs(19) <= '0';
            xs(20) <= '0';   

        when "0011"&"0101" => --t5q3
            xs(0)  <= '0';
            xs(1)  <= '0';
            xs(2)  <= '0';
            xs(3)  <= '0';
            xs(4)  <= '0';
            xs(5)  <= '0';
            xs(6)  <= '0';
            xs(7)  <= '0';
            xs(8)  <= '0';
            xs(9)  <= '0';
            xs(10) <= '1';
            xs(11) <= '0';
            xs(12) <= '0';
            xs(13) <= '0';
            xs(14) <= '0';
            xs(15) <= '0';
            xs(16) <= '0';
            xs(17) <= '0';
            xs(18) <= '0';
            xs(19) <= '0';
            xs(20) <= '0'; 
            
        when "0011"&"0110" => --t6q3
            xs(0)  <= '0';
            xs(1)  <= '0';
            xs(2)  <= '0';
            xs(3)  <= '0';
            xs(4)  <= '0';
            xs(5)  <= '0';
            xs(6)  <= '0';
            xs(7)  <= '0';
            xs(8)  <= '1';
            xs(9)  <= '0';
            xs(10) <= '0';
            xs(11) <= '0';
            xs(12) <= '0';
            xs(13) <= '0';
            xs(14) <= '0';
            xs(15) <= '0';
            xs(16) <= '0';
            xs(17) <= '0';
            xs(18) <= '0';
            xs(19) <= '0';
            xs(20) <= '0'; 
            
        when "0011"&"0111" => --t7q3
            xs(0)  <= '0';
            xs(1)  <= '0';
            xs(2)  <= '1';
            xs(3)  <= '0';
            xs(4)  <= '0';
            xs(5)  <= '0';
            xs(6)  <= '1';
            xs(7)  <= '0';
            xs(8)  <= '0';
            xs(9)  <= '0';
            xs(10) <= '0';
            xs(11) <= '0';
            xs(12) <= '0';
            xs(13) <= '0';
            xs(14) <= '0';
            xs(15) <= '0';
            xs(16) <= '0';
            xs(17) <= '0';
            xs(18) <= '0';
            xs(19) <= '0';
            xs(20) <= '0'; 

        when "0011"&"1000" => --t8q3
            xs(0)  <= '0';
            xs(1)  <= '0';
            xs(2)  <= '0';
            xs(3)  <= '0';
            xs(4)  <= '0';
            xs(5)  <= '0';
            xs(6)  <= '0';
            xs(7)  <= '1';
            xs(8)  <= '0';
            xs(9)  <= '0';
            xs(10) <= '0';
            xs(11) <= '0';
            xs(12) <= '0';
            xs(13) <= '0';
            xs(14) <= '0';
            xs(15) <= '0';
            xs(16) <= '0';
            xs(17) <= '0';
            xs(18) <= '0';
            xs(19) <= '0';
            xs(20) <= '0'; 

        when "0011"&"1001" => --t9q3
            xs(0)  <= '0';
            xs(1)  <= '1';
            xs(2)  <= '0';
            xs(3)  <= '0';
            xs(4)  <= '0';
            xs(5)  <= '0';
            xs(6)  <= '0';
            xs(7)  <= '0';
            xs(8)  <= '0';
            xs(9)  <= '0';
            xs(10) <= '0';
            xs(11) <= '0';
            xs(12) <= '0';
            xs(13) <= '0';
            xs(14) <= '0';
            xs(15) <= '0';
            xs(16) <= '0';
            xs(17) <= '0';
            xs(18) <= '0';
            xs(19) <= '0';
            xs(20) <= '0'; 

        when "0011"&"1010" => --tAq3
            xs(0)  <= '0';
            xs(1)  <= '0';
            xs(2)  <= '0';
            xs(3)  <= '0';
            xs(4)  <= '0';
            xs(5)  <= '0';
            xs(6)  <= '0';
            xs(7)  <= '0';
            xs(8)  <= '0';
            xs(9)  <= '0';
            xs(10) <= '0';
            xs(11) <= '0';
            xs(12) <= '0';
            xs(13) <= '0';
            xs(14) <= '0';
            xs(15) <= '0';
            xs(16) <= '0';
            xs(17) <= '0';
            xs(18) <= '0';
            xs(19) <= '0';
            xs(20) <= '1'; 

        when "0011"&"1011" => --tBq3
            xs(0)  <= '0';
            xs(1)  <= '0';
            xs(2)  <= '0';
            xs(3)  <= '0';
            xs(4)  <= '0';
            xs(5)  <= '0';
            xs(6)  <= '0';
            xs(7)  <= '0';
            xs(8)  <= '0';
            xs(9)  <= '0';
            xs(10) <= '0';
            xs(11) <= '0';
            xs(12) <= '0';
            xs(13) <= '0';
            xs(14) <= '1';
            xs(15) <= '0';
            xs(16) <= '0';
            xs(17) <= '0';
            xs(18) <= '0';
            xs(19) <= '0';
            xs(20) <= '0'; 
------------  FIN -> 03h  MOV [DIR], A            
            
------------ 04h  XOR A, N     
        --       q & t
        when "0100"&"0000" => --t0
            xs(0)  <= '0';
            xs(1)  <= '0';
            xs(2)  <= '0';
            xs(3)  <= '0';
            xs(4)  <= '0';
            xs(5)  <= '0';
            xs(6)  <= '0';
            xs(7)  <= '0';
            xs(8)  <= '1';
            xs(9)  <= '0';
            xs(10) <= '0';
            xs(11) <= '0';
            xs(12) <= '0';
            xs(13) <= '0';
            xs(14) <= '0';
            xs(15) <= '0';
            xs(16) <= '0';
            xs(17) <= '0';
            xs(18) <= '0';
            xs(19) <= '0';
            xs(20) <= '0';

        when "0100"&"0001" => --t1
            xs(0)  <= '0';
            xs(1)  <= '0';
            xs(2)  <= '1';
            xs(3)  <= '0';
            xs(4)  <= '0';
            xs(5)  <= '0';
            xs(6)  <= '1';
            xs(7)  <= '0';
            xs(8)  <= '0';
            xs(9)  <= '0';
            xs(10) <= '0';
            xs(11) <= '0';
            xs(12) <= '0';
            xs(13) <= '0';
            xs(14) <= '0';
            xs(15) <= '0';
            xs(16) <= '0';
            xs(17) <= '0';
            xs(18) <= '0';
            xs(19) <= '0';
            xs(20) <= '0';    
            
        when "0100"&"0010" => --t2
            xs(0)  <= '1';
            xs(1)  <= '0';
            xs(2)  <= '0';
            xs(3)  <= '0';
            xs(4)  <= '0';
            xs(5)  <= '0';
            xs(6)  <= '0';
            xs(7)  <= '0';
            xs(8)  <= '0';
            xs(9)  <= '0';
            xs(10) <= '0';
            xs(11) <= '0';
            xs(12) <= '0';
            xs(13) <= '0';
            xs(14) <= '0';
            xs(15) <= '0';
            xs(16) <= '0';
            xs(17) <= '0';
            xs(18) <= '0';
            xs(19) <= '0';
            xs(20) <= '0';    
            
        when "0100"&"0011" => --t3q4
            xs(0)  <= '0';
            xs(1)  <= '0';
            xs(2)  <= '0';
            xs(3)  <= '0';
            xs(4)  <= '0';
            xs(5)  <= '0';
            xs(6)  <= '0';
            xs(7)  <= '0';
            xs(8)  <= '1';
            xs(9)  <= '0';
            xs(10) <= '0';
            xs(11) <= '0';
            xs(12) <= '0';
            xs(13) <= '0';
            xs(14) <= '0';
            xs(15) <= '0';
            xs(16) <= '0';
            xs(17) <= '0';
            xs(18) <= '0';
            xs(19) <= '0';
            xs(20) <= '0';  
            
        when "0100"&"0100" => --t4q4
            xs(0)  <= '0';
            xs(1)  <= '0';
            xs(2)  <= '1';
            xs(3)  <= '0';
            xs(4)  <= '0';
            xs(5)  <= '0';
            xs(6)  <= '1';
            xs(7)  <= '0';
            xs(8)  <= '0';
            xs(9)  <= '0';
            xs(10) <= '0';
            xs(11) <= '0';
            xs(12) <= '0';
            xs(13) <= '0';
            xs(14) <= '0';
            xs(15) <= '0';
            xs(16) <= '0';
            xs(17) <= '0';
            xs(18) <= '0';
            xs(19) <= '0';
            xs(20) <= '0';   

        when "0100"&"0101" => --t5q4
            xs(0)  <= '0';
            xs(1)  <= '0';
            xs(2)  <= '0';
            xs(3)  <= '0';
            xs(4)  <= '0';
            xs(5)  <= '0';
            xs(6)  <= '0';
            xs(7)  <= '0';
            xs(8)  <= '0';
            xs(9)  <= '0';
            xs(10) <= '0';
            xs(11) <= '0';
            xs(12) <= '0';
            xs(13) <= '0';
            xs(14) <= '0';
            xs(15) <= '1';
            xs(16) <= '1';
            xs(17) <= '0';
            xs(18) <= '0';
            xs(19) <= '1';
            xs(20) <= '0'; 
            
        when "0100"&"0110" => --t6q4
            xs(0)  <= '0';
            xs(1)  <= '0';
            xs(2)  <= '0';
            xs(3)  <= '0';
            xs(4)  <= '0';
            xs(5)  <= '0';
            xs(6)  <= '0';
            xs(7)  <= '0';
            xs(8)  <= '0';
            xs(9)  <= '0';
            xs(10) <= '0';
            xs(11) <= '0';
            xs(12) <= '0';
            xs(13) <= '0';
            xs(14) <= '1';
            xs(15) <= '0';
            xs(16) <= '0';
            xs(17) <= '0';
            xs(18) <= '0';
            xs(19) <= '0';
            xs(20) <= '0'; 
------------  FIN -> 04h  XOR A, N        
            
------------ 05h  ADD A, [DIR]    
        --       q & t
        when "0101"&"0000" => --t0
            xs(0)  <= '0';
            xs(1)  <= '0';
            xs(2)  <= '0';
            xs(3)  <= '0';
            xs(4)  <= '0';
            xs(5)  <= '0';
            xs(6)  <= '0';
            xs(7)  <= '0';
            xs(8)  <= '1';
            xs(9)  <= '0';
            xs(10) <= '0';
            xs(11) <= '0';
            xs(12) <= '0';
            xs(13) <= '0';
            xs(14) <= '0';
            xs(15) <= '0';
            xs(16) <= '0';
            xs(17) <= '0';
            xs(18) <= '0';
            xs(19) <= '0';
            xs(20) <= '0';

        when "0101"&"0001" => --t1
            xs(0)  <= '0';
            xs(1)  <= '0';
            xs(2)  <= '1';
            xs(3)  <= '0';
            xs(4)  <= '0';
            xs(5)  <= '0';
            xs(6)  <= '1';
            xs(7)  <= '0';
            xs(8)  <= '0';
            xs(9)  <= '0';
            xs(10) <= '0';
            xs(11) <= '0';
            xs(12) <= '0';
            xs(13) <= '0';
            xs(14) <= '0';
            xs(15) <= '0';
            xs(16) <= '0';
            xs(17) <= '0';
            xs(18) <= '0';
            xs(19) <= '0';
            xs(20) <= '0';    
            
        when "0101"&"0010" => --t2
            xs(0)  <= '1';
            xs(1)  <= '0';
            xs(2)  <= '0';
            xs(3)  <= '0';
            xs(4)  <= '0';
            xs(5)  <= '0';
            xs(6)  <= '0';
            xs(7)  <= '0';
            xs(8)  <= '0';
            xs(9)  <= '0';
            xs(10) <= '0';
            xs(11) <= '0';
            xs(12) <= '0';
            xs(13) <= '0';
            xs(14) <= '0';
            xs(15) <= '0';
            xs(16) <= '0';
            xs(17) <= '0';
            xs(18) <= '0';
            xs(19) <= '0';
            xs(20) <= '0';    
            
        when "0101"&"0011" => --t3q5
            xs(0)  <= '0';
            xs(1)  <= '0';
            xs(2)  <= '0';
            xs(3)  <= '0';
            xs(4)  <= '0';
            xs(5)  <= '0';
            xs(6)  <= '0';
            xs(7)  <= '0';
            xs(8)  <= '1';
            xs(9)  <= '0';
            xs(10) <= '0';
            xs(11) <= '0';
            xs(12) <= '0';
            xs(13) <= '0';
            xs(14) <= '0';
            xs(15) <= '0';
            xs(16) <= '0';
            xs(17) <= '0';
            xs(18) <= '0';
            xs(19) <= '0';
            xs(20) <= '0';  
            
        when "0101"&"0100" => --t4q5
            xs(0)  <= '0';
            xs(1)  <= '0';
            xs(2)  <= '1';
            xs(3)  <= '0';
            xs(4)  <= '0';
            xs(5)  <= '0';
            xs(6)  <= '1';
            xs(7)  <= '0';
            xs(8)  <= '0';
            xs(9)  <= '0';
            xs(10) <= '0';
            xs(11) <= '0';
            xs(12) <= '0';
            xs(13) <= '0';
            xs(14) <= '0';
            xs(15) <= '0';
            xs(16) <= '0';
            xs(17) <= '0';
            xs(18) <= '0';
            xs(19) <= '0';
            xs(20) <= '0';   

        when "0101"&"0101" => --t5q5
            xs(0)  <= '0';
            xs(1)  <= '0';
            xs(2)  <= '0';
            xs(3)  <= '0';
            xs(4)  <= '0';
            xs(5)  <= '0';
            xs(6)  <= '0';
            xs(7)  <= '0';
            xs(8)  <= '0';
            xs(9)  <= '0';
            xs(10) <= '1';
            xs(11) <= '0';
            xs(12) <= '0';
            xs(13) <= '0';
            xs(14) <= '0';
            xs(15) <= '0';
            xs(16) <= '0';
            xs(17) <= '0';
            xs(18) <= '0';
            xs(19) <= '0';
            xs(20) <= '0'; 
            
        when "0101"&"0110" => --t6q5
            xs(0)  <= '0';
            xs(1)  <= '0';
            xs(2)  <= '0';
            xs(3)  <= '0';
            xs(4)  <= '0';
            xs(5)  <= '0';
            xs(6)  <= '0';
            xs(7)  <= '0';
            xs(8)  <= '1';
            xs(9)  <= '0';
            xs(10) <= '0';
            xs(11) <= '0';
            xs(12) <= '0';
            xs(13) <= '0';
            xs(14) <= '0';
            xs(15) <= '0';
            xs(16) <= '0';
            xs(17) <= '0';
            xs(18) <= '0';
            xs(19) <= '0';
            xs(20) <= '0'; 

        when "0101"&"0111" => --t7q5
            xs(0)  <= '0';
            xs(1)  <= '0';
            xs(2)  <= '1';
            xs(3)  <= '0';
            xs(4)  <= '0';
            xs(5)  <= '0';
            xs(6)  <= '1';
            xs(7)  <= '0';
            xs(8)  <= '0';
            xs(9)  <= '0';
            xs(10) <= '0';
            xs(11) <= '0';
            xs(12) <= '0';
            xs(13) <= '0';
            xs(14) <= '0';
            xs(15) <= '0';
            xs(16) <= '0';
            xs(17) <= '0';
            xs(18) <= '0';
            xs(19) <= '0';
            xs(20) <= '0'; 

        when "0101"&"1000" => --t8q5
            xs(0)  <= '0';
            xs(1)  <= '0';
            xs(2)  <= '0';
            xs(3)  <= '0';
            xs(4)  <= '0';
            xs(5)  <= '0';
            xs(6)  <= '0';
            xs(7)  <= '1';
            xs(8)  <= '0';
            xs(9)  <= '0';
            xs(10) <= '0';
            xs(11) <= '0';
            xs(12) <= '0';
            xs(13) <= '0';
            xs(14) <= '0';
            xs(15) <= '0';
            xs(16) <= '0';
            xs(17) <= '0';
            xs(18) <= '0';
            xs(19) <= '0';
            xs(20) <= '0'; 

        when "0101"&"1001" => --t9q5
            xs(0)  <= '0';
            xs(1)  <= '0';
            xs(2)  <= '1';
            xs(3)  <= '0';
            xs(4)  <= '0';
            xs(5)  <= '0';
            xs(6)  <= '0';
            xs(7)  <= '0';
            xs(8)  <= '0';
            xs(9)  <= '0';
            xs(10) <= '0';
            xs(11) <= '0';
            xs(12) <= '0';
            xs(13) <= '0';
            xs(14) <= '0';
            xs(15) <= '0';
            xs(16) <= '0';
            xs(17) <= '0';
            xs(18) <= '0';
            xs(19) <= '0';
            xs(20) <= '0'; 

        when "0101"&"1010" => --tAq5
            xs(0)  <= '0';
            xs(1)  <= '0';
            xs(2)  <= '0';
            xs(3)  <= '0';
            xs(4)  <= '0';
            xs(5)  <= '0';
            xs(6)  <= '0';
            xs(7)  <= '0';
            xs(8)  <= '0';
            xs(9)  <= '0';
            xs(10) <= '0';
            xs(11) <= '0';
            xs(12) <= '0';
            xs(13) <= '0';
            xs(14) <= '0';
            xs(15) <= '0';
            xs(16) <= '1';
            xs(17) <= '1';
            xs(18) <= '0';
            xs(19) <= '1';
            xs(20) <= '0'; 

        when "0101"&"1011" => --tBq5
            xs(0)  <= '0';
            xs(1)  <= '0';
            xs(2)  <= '0';
            xs(3)  <= '0';
            xs(4)  <= '0';
            xs(5)  <= '0';
            xs(6)  <= '0';
            xs(7)  <= '0';
            xs(8)  <= '0';
            xs(9)  <= '0';
            xs(10) <= '0';
            xs(11) <= '0';
            xs(12) <= '0';
            xs(13) <= '0';
            xs(14) <= '1';
            xs(15) <= '0';
            xs(16) <= '0';
            xs(17) <= '0';
            xs(18) <= '0';
            xs(19) <= '0';
            xs(20) <= '0'; 
------------  FIN -> 05h  ADD A, [DIR]   
    
------------ 06h  AND A, [DIR]    
        --       q & t
        when "0110"&"0000" => --t0
            xs(0)  <= '0';
            xs(1)  <= '0';
            xs(2)  <= '0';
            xs(3)  <= '0';
            xs(4)  <= '0';
            xs(5)  <= '0';
            xs(6)  <= '0';
            xs(7)  <= '0';
            xs(8)  <= '1';
            xs(9)  <= '0';
            xs(10) <= '0';
            xs(11) <= '0';
            xs(12) <= '0';
            xs(13) <= '0';
            xs(14) <= '0';
            xs(15) <= '0';
            xs(16) <= '0';
            xs(17) <= '0';
            xs(18) <= '0';
            xs(19) <= '0';
            xs(20) <= '0';

        when "0110"&"0001" => --t1
            xs(0)  <= '0';
            xs(1)  <= '0';
            xs(2)  <= '1';
            xs(3)  <= '0';
            xs(4)  <= '0';
            xs(5)  <= '0';
            xs(6)  <= '1';
            xs(7)  <= '0';
            xs(8)  <= '0';
            xs(9)  <= '0';
            xs(10) <= '0';
            xs(11) <= '0';
            xs(12) <= '0';
            xs(13) <= '0';
            xs(14) <= '0';
            xs(15) <= '0';
            xs(16) <= '0';
            xs(17) <= '0';
            xs(18) <= '0';
            xs(19) <= '0';
            xs(20) <= '0';    
            
        when "0110"&"0010" => --t2
            xs(0)  <= '1';
            xs(1)  <= '0';
            xs(2)  <= '0';
            xs(3)  <= '0';
            xs(4)  <= '0';
            xs(5)  <= '0';
            xs(6)  <= '0';
            xs(7)  <= '0';
            xs(8)  <= '0';
            xs(9)  <= '0';
            xs(10) <= '0';
            xs(11) <= '0';
            xs(12) <= '0';
            xs(13) <= '0';
            xs(14) <= '0';
            xs(15) <= '0';
            xs(16) <= '0';
            xs(17) <= '0';
            xs(18) <= '0';
            xs(19) <= '0';
            xs(20) <= '0';    
            
        when "0110"&"0011" => --t3q6
            xs(0)  <= '0';
            xs(1)  <= '0';
            xs(2)  <= '1';
            xs(3)  <= '0';
            xs(4)  <= '0';
            xs(5)  <= '0';
            xs(6)  <= '1';
            xs(7)  <= '0';
            xs(8)  <= '0';
            xs(9)  <= '0';
            xs(10) <= '0';
            xs(11) <= '0';
            xs(12) <= '0';
            xs(13) <= '0';
            xs(14) <= '0';
            xs(15) <= '0';
            xs(16) <= '0';
            xs(17) <= '0';
            xs(18) <= '0';
            xs(19) <= '0';
            xs(20) <= '0';  
            
        when "0110"&"0100" => --t4q6
            xs(0)  <= '0';
            xs(1)  <= '0';
            xs(2)  <= '1';
            xs(3)  <= '0';
            xs(4)  <= '0';
            xs(5)  <= '0';
            xs(6)  <= '1';
            xs(7)  <= '0';
            xs(8)  <= '0';
            xs(9)  <= '0';
            xs(10) <= '0';
            xs(11) <= '0';
            xs(12) <= '0';
            xs(13) <= '0';
            xs(14) <= '0';
            xs(15) <= '0';
            xs(16) <= '0';
            xs(17) <= '0';
            xs(18) <= '0';
            xs(19) <= '0';
            xs(20) <= '0';   

        when "0110"&"0101" => --t5q6
            xs(0)  <= '0';
            xs(1)  <= '0';
            xs(2)  <= '0';
            xs(3)  <= '0';
            xs(4)  <= '0';
            xs(5)  <= '0';
            xs(6)  <= '0';
            xs(7)  <= '0';
            xs(8)  <= '0';
            xs(9)  <= '0';
            xs(10) <= '1';
            xs(11) <= '0';
            xs(12) <= '0';
            xs(13) <= '0';
            xs(14) <= '0';
            xs(15) <= '0';
            xs(16) <= '0';
            xs(17) <= '0';
            xs(18) <= '0';
            xs(19) <= '0';
            xs(20) <= '0'; 
            
        when "0110"&"0110" => --t6q6
            xs(0)  <= '0';
            xs(1)  <= '0';
            xs(2)  <= '0';
            xs(3)  <= '0';
            xs(4)  <= '0';
            xs(5)  <= '0';
            xs(6)  <= '0';
            xs(7)  <= '0';
            xs(8)  <= '1';
            xs(9)  <= '0';
            xs(10) <= '0';
            xs(11) <= '0';
            xs(12) <= '0';
            xs(13) <= '0';
            xs(14) <= '0';
            xs(15) <= '0';
            xs(16) <= '0';
            xs(17) <= '0';
            xs(18) <= '0';
            xs(19) <= '0';
            xs(20) <= '0'; 

        when "0110"&"0111" => --t7q6
            xs(0)  <= '0';
            xs(1)  <= '0';
            xs(2)  <= '1';
            xs(3)  <= '0';
            xs(4)  <= '0';
            xs(5)  <= '0';
            xs(6)  <= '1';
            xs(7)  <= '0';
            xs(8)  <= '0';
            xs(9)  <= '0';
            xs(10) <= '0';
            xs(11) <= '0';
            xs(12) <= '0';
            xs(13) <= '0';
            xs(14) <= '0';
            xs(15) <= '0';
            xs(16) <= '0';
            xs(17) <= '0';
            xs(18) <= '0';
            xs(19) <= '0';
            xs(20) <= '0'; 

        when "0110"&"1000" => --t8q6
            xs(0)  <= '0';
            xs(1)  <= '0';
            xs(2)  <= '0';
            xs(3)  <= '0';
            xs(4)  <= '0';
            xs(5)  <= '0';
            xs(6)  <= '0';
            xs(7)  <= '1';
            xs(8)  <= '0';
            xs(9)  <= '0';
            xs(10) <= '0';
            xs(11) <= '0';
            xs(12) <= '0';
            xs(13) <= '0';
            xs(14) <= '0';
            xs(15) <= '0';
            xs(16) <= '0';
            xs(17) <= '0';
            xs(18) <= '0';
            xs(19) <= '0';
            xs(20) <= '0'; 

        when "0110"&"1001" => --t9q6
            xs(0)  <= '0';
            xs(1)  <= '0';
            xs(2)  <= '1';
            xs(3)  <= '0';
            xs(4)  <= '0';
            xs(5)  <= '0';
            xs(6)  <= '0';
            xs(7)  <= '0';
            xs(8)  <= '0';
            xs(9)  <= '0';
            xs(10) <= '0';
            xs(11) <= '0';
            xs(12) <= '0';
            xs(13) <= '0';
            xs(14) <= '0';
            xs(15) <= '0';
            xs(16) <= '0';
            xs(17) <= '0';
            xs(18) <= '0';
            xs(19) <= '0';
            xs(20) <= '0'; 

        when "0110"&"1010" => --tAq6
            xs(0)  <= '0';
            xs(1)  <= '0';
            xs(2)  <= '0';
            xs(3)  <= '0';
            xs(4)  <= '0';
            xs(5)  <= '0';
            xs(6)  <= '0';
            xs(7)  <= '0';
            xs(8)  <= '0';
            xs(9)  <= '0';
            xs(10) <= '0';
            xs(11) <= '0';
            xs(12) <= '0';
            xs(13) <= '0';
            xs(14) <= '0';
            xs(15) <= '1';
            xs(16) <= '0';
            xs(17) <= '0';
            xs(18) <= '0';
            xs(19) <= '1';
            xs(20) <= '0'; 

        when "0110"&"1011" => --tBq6
            xs(0)  <= '0';
            xs(1)  <= '0';
            xs(2)  <= '0';
            xs(3)  <= '0';
            xs(4)  <= '0';
            xs(5)  <= '0';
            xs(6)  <= '0';
            xs(7)  <= '0';
            xs(8)  <= '0';
            xs(9)  <= '0';
            xs(10) <= '0';
            xs(11) <= '0';
            xs(12) <= '0';
            xs(13) <= '0';
            xs(14) <= '1';
            xs(15) <= '0';
            xs(16) <= '0';
            xs(17) <= '0';
            xs(18) <= '0';
            xs(19) <= '0';
            xs(20) <= '0'; 
------------  FIN -> 06h  AND A, [DIR]  

------------ 07h  OR A, [DIR]   
        --       q & t
        when "0111"&"0000" => --t0
            xs(0)  <= '0';
            xs(1)  <= '0';
            xs(2)  <= '0';
            xs(3)  <= '0';
            xs(4)  <= '0';
            xs(5)  <= '0';
            xs(6)  <= '0';
            xs(7)  <= '0';
            xs(8)  <= '1';
            xs(9)  <= '0';
            xs(10) <= '0';
            xs(11) <= '0';
            xs(12) <= '0';
            xs(13) <= '0';
            xs(14) <= '0';
            xs(15) <= '0';
            xs(16) <= '0';
            xs(17) <= '0';
            xs(18) <= '0';
            xs(19) <= '0';
            xs(20) <= '0';

        when "0111"&"0001" => --t1
            xs(0)  <= '0';
            xs(1)  <= '0';
            xs(2)  <= '1';
            xs(3)  <= '0';
            xs(4)  <= '0';
            xs(5)  <= '0';
            xs(6)  <= '1';
            xs(7)  <= '0';
            xs(8)  <= '0';
            xs(9)  <= '0';
            xs(10) <= '0';
            xs(11) <= '0';
            xs(12) <= '0';
            xs(13) <= '0';
            xs(14) <= '0';
            xs(15) <= '0';
            xs(16) <= '0';
            xs(17) <= '0';
            xs(18) <= '0';
            xs(19) <= '0';
            xs(20) <= '0';    
            
        when "0111"&"0010" => --t2
            xs(0)  <= '1';
            xs(1)  <= '0';
            xs(2)  <= '0';
            xs(3)  <= '0';
            xs(4)  <= '0';
            xs(5)  <= '0';
            xs(6)  <= '0';
            xs(7)  <= '0';
            xs(8)  <= '0';
            xs(9)  <= '0';
            xs(10) <= '0';
            xs(11) <= '0';
            xs(12) <= '0';
            xs(13) <= '0';
            xs(14) <= '0';
            xs(15) <= '0';
            xs(16) <= '0';
            xs(17) <= '0';
            xs(18) <= '0';
            xs(19) <= '0';
            xs(20) <= '0';    
            
        when "0111"&"0011" => --t3q7
            xs(0)  <= '0';
            xs(1)  <= '0';
            xs(2)  <= '0';
            xs(3)  <= '0';
            xs(4)  <= '0';
            xs(5)  <= '0';
            xs(6)  <= '0';
            xs(7)  <= '0';
            xs(8)  <= '1';
            xs(9)  <= '0';
            xs(10) <= '0';
            xs(11) <= '0';
            xs(12) <= '0';
            xs(13) <= '0';
            xs(14) <= '0';
            xs(15) <= '0';
            xs(16) <= '0';
            xs(17) <= '0';
            xs(18) <= '0';
            xs(19) <= '0';
            xs(20) <= '0';  
            
        when "0111"&"0100" => --t4q7
            xs(0)  <= '0';
            xs(1)  <= '0';
            xs(2)  <= '1';
            xs(3)  <= '0';
            xs(4)  <= '0';
            xs(5)  <= '0';
            xs(6)  <= '1';
            xs(7)  <= '0';
            xs(8)  <= '0';
            xs(9)  <= '0';
            xs(10) <= '0';
            xs(11) <= '0';
            xs(12) <= '0';
            xs(13) <= '0';
            xs(14) <= '0';
            xs(15) <= '0';
            xs(16) <= '0';
            xs(17) <= '0';
            xs(18) <= '0';
            xs(19) <= '0';
            xs(20) <= '0';   

        when "0111"&"0101" => --t5q7
            xs(0)  <= '0';
            xs(1)  <= '0';
            xs(2)  <= '0';
            xs(3)  <= '0';
            xs(4)  <= '0';
            xs(5)  <= '0';
            xs(6)  <= '0';
            xs(7)  <= '0';
            xs(8)  <= '0';
            xs(9)  <= '0';
            xs(10) <= '1';
            xs(11) <= '0';
            xs(12) <= '0';
            xs(13) <= '0';
            xs(14) <= '0';
            xs(15) <= '0';
            xs(16) <= '0';
            xs(17) <= '0';
            xs(18) <= '0';
            xs(19) <= '0';
            xs(20) <= '0'; 
            
        when "0111"&"0110" => --t6q7
            xs(0)  <= '0';
            xs(1)  <= '0';
            xs(2)  <= '0';
            xs(3)  <= '0';
            xs(4)  <= '0';
            xs(5)  <= '0';
            xs(6)  <= '0';
            xs(7)  <= '0';
            xs(8)  <= '1';
            xs(9)  <= '0';
            xs(10) <= '0';
            xs(11) <= '0';
            xs(12) <= '0';
            xs(13) <= '0';
            xs(14) <= '0';
            xs(15) <= '0';
            xs(16) <= '0';
            xs(17) <= '0';
            xs(18) <= '0';
            xs(19) <= '0';
            xs(20) <= '0'; 

        when "0111"&"0111" => --t7q7
            xs(0)  <= '0';
            xs(1)  <= '0';
            xs(2)  <= '1';
            xs(3)  <= '0';
            xs(4)  <= '0';
            xs(5)  <= '0';
            xs(6)  <= '1';
            xs(7)  <= '0';
            xs(8)  <= '0';
            xs(9)  <= '0';
            xs(10) <= '0';
            xs(11) <= '0';
            xs(12) <= '0';
            xs(13) <= '0';
            xs(14) <= '0';
            xs(15) <= '0';
            xs(16) <= '0';
            xs(17) <= '0';
            xs(18) <= '0';
            xs(19) <= '0';
            xs(20) <= '0'; 

        when "0111"&"1000" => --t8q7
            xs(0)  <= '0';
            xs(1)  <= '0';
            xs(2)  <= '0';
            xs(3)  <= '0';
            xs(4)  <= '0';
            xs(5)  <= '0';
            xs(6)  <= '0';
            xs(7)  <= '1';
            xs(8)  <= '0';
            xs(9)  <= '0';
            xs(10) <= '0';
            xs(11) <= '0';
            xs(12) <= '0';
            xs(13) <= '0';
            xs(14) <= '0';
            xs(15) <= '0';
            xs(16) <= '0';
            xs(17) <= '0';
            xs(18) <= '0';
            xs(19) <= '0';
            xs(20) <= '0'; 

        when "0111"&"1001" => --t9q7
            xs(0)  <= '0';
            xs(1)  <= '0';
            xs(2)  <= '1';
            xs(3)  <= '0';
            xs(4)  <= '0';
            xs(5)  <= '0';
            xs(6)  <= '0';
            xs(7)  <= '0';
            xs(8)  <= '0';
            xs(9)  <= '0';
            xs(10) <= '0';
            xs(11) <= '0';
            xs(12) <= '0';
            xs(13) <= '0';
            xs(14) <= '0';
            xs(15) <= '0';
            xs(16) <= '0';
            xs(17) <= '0';
            xs(18) <= '0';
            xs(19) <= '0';
            xs(20) <= '0'; 

        when "0111"&"1010" => --tAq7
            xs(0)  <= '0';
            xs(1)  <= '0';
            xs(2)  <= '0';
            xs(3)  <= '0';
            xs(4)  <= '0';
            xs(5)  <= '0';
            xs(6)  <= '0';
            xs(7)  <= '0';
            xs(8)  <= '0';
            xs(9)  <= '0';
            xs(10) <= '0';
            xs(11) <= '0';
            xs(12) <= '0';
            xs(13) <= '0';
            xs(14) <= '0';
            xs(15) <= '0';
            xs(16) <= '1';
            xs(17) <= '0';
            xs(18) <= '0';
            xs(19) <= '1';
            xs(20) <= '0'; 

        when "0111"&"1011" => --tBq7
            xs(0)  <= '0';
            xs(1)  <= '0';
            xs(2)  <= '0';
            xs(3)  <= '0';
            xs(4)  <= '0';
            xs(5)  <= '0';
            xs(6)  <= '0';
            xs(7)  <= '0';
            xs(8)  <= '0';
            xs(9)  <= '0';
            xs(10) <= '0';
            xs(11) <= '0';
            xs(12) <= '0';
            xs(13) <= '0';
            xs(14) <= '1';
            xs(15) <= '0';
            xs(16) <= '0';
            xs(17) <= '0';
            xs(18) <= '0';
            xs(19) <= '0';
            xs(20) <= '0'; 
------------  FIN -> 07h  OR A, [DIR]  

------------ 08h  JMP DIR   
        --       q & t
        when "1000"&"0000" => --t0
            xs(0)  <= '0';
            xs(1)  <= '0';
            xs(2)  <= '0';
            xs(3)  <= '0';
            xs(4)  <= '0';
            xs(5)  <= '0';
            xs(6)  <= '0';
            xs(7)  <= '0';
            xs(8)  <= '1';
            xs(9)  <= '0';
            xs(10) <= '0';
            xs(11) <= '0';
            xs(12) <= '0';
            xs(13) <= '0';
            xs(14) <= '0';
            xs(15) <= '0';
            xs(16) <= '0';
            xs(17) <= '0';
            xs(18) <= '0';
            xs(19) <= '0';
            xs(20) <= '0';

        when "1000"&"0001" => --t1
            xs(0)  <= '0';
            xs(1)  <= '0';
            xs(2)  <= '1';
            xs(3)  <= '0';
            xs(4)  <= '0';
            xs(5)  <= '0';
            xs(6)  <= '1';
            xs(7)  <= '0';
            xs(8)  <= '0';
            xs(9)  <= '0';
            xs(10) <= '0';
            xs(11) <= '0';
            xs(12) <= '0';
            xs(13) <= '0';
            xs(14) <= '0';
            xs(15) <= '0';
            xs(16) <= '0';
            xs(17) <= '0';
            xs(18) <= '0';
            xs(19) <= '0';
            xs(20) <= '0';    
            
        when "1000"&"0010" => --t2
            xs(0)  <= '1';
            xs(1)  <= '0';
            xs(2)  <= '0';
            xs(3)  <= '0';
            xs(4)  <= '0';
            xs(5)  <= '0';
            xs(6)  <= '0';
            xs(7)  <= '0';
            xs(8)  <= '0';
            xs(9)  <= '0';
            xs(10) <= '0';
            xs(11) <= '0';
            xs(12) <= '0';
            xs(13) <= '0';
            xs(14) <= '0';
            xs(15) <= '0';
            xs(16) <= '0';
            xs(17) <= '0';
            xs(18) <= '0';
            xs(19) <= '0';
            xs(20) <= '0';    
            
        when "1000"&"0011" => --t3q8
            xs(0)  <= '0';
            xs(1)  <= '0';
            xs(2)  <= '0';
            xs(3)  <= '0';
            xs(4)  <= '0';
            xs(5)  <= '0';
            xs(6)  <= '0';
            xs(7)  <= '0';
            xs(8)  <= '1';
            xs(9)  <= '0';
            xs(10) <= '0';
            xs(11) <= '0';
            xs(12) <= '0';
            xs(13) <= '0';
            xs(14) <= '0';
            xs(15) <= '0';
            xs(16) <= '0';
            xs(17) <= '0';
            xs(18) <= '0';
            xs(19) <= '0';
            xs(20) <= '0';  
            
        when "1000"&"0100" => --t4q8
            xs(0)  <= '0';
            xs(1)  <= '0';
            xs(2)  <= '1';
            xs(3)  <= '0';
            xs(4)  <= '0';
            xs(5)  <= '0';
            xs(6)  <= '1';
            xs(7)  <= '0';
            xs(8)  <= '0';
            xs(9)  <= '0';
            xs(10) <= '0';
            xs(11) <= '0';
            xs(12) <= '0';
            xs(13) <= '0';
            xs(14) <= '0';
            xs(15) <= '0';
            xs(16) <= '0';
            xs(17) <= '0';
            xs(18) <= '0';
            xs(19) <= '0';
            xs(20) <= '0';   

        when "1000"&"0101" => --t5q8
            xs(0)  <= '0';
            xs(1)  <= '0';
            xs(2)  <= '0';
            xs(3)  <= '0';
            xs(4)  <= '0';
            xs(5)  <= '0';
            xs(6)  <= '0';
            xs(7)  <= '0';
            xs(8)  <= '0';
            xs(9)  <= '0';
            xs(10) <= '1';
            xs(11) <= '0';
            xs(12) <= '0';
            xs(13) <= '0';
            xs(14) <= '0';
            xs(15) <= '0';
            xs(16) <= '0';
            xs(17) <= '0';
            xs(18) <= '0';
            xs(19) <= '0';
            xs(20) <= '0'; 
            
        when "1000"&"0110" => --t6q8
            xs(0)  <= '0';
            xs(1)  <= '0';
            xs(2)  <= '0';
            xs(3)  <= '0';
            xs(4)  <= '0';
            xs(5)  <= '0';
            xs(6)  <= '0';
            xs(7)  <= '0';
            xs(8)  <= '1';
            xs(9)  <= '0';
            xs(10) <= '0';
            xs(11) <= '0';
            xs(12) <= '0';
            xs(13) <= '0';
            xs(14) <= '0';
            xs(15) <= '0';
            xs(16) <= '0';
            xs(17) <= '0';
            xs(18) <= '0';
            xs(19) <= '0';
            xs(20) <= '0'; 

        when "1000"&"0111" => --t7q8
            xs(0)  <= '0';
            xs(1)  <= '0';
            xs(2)  <= '1';
            xs(3)  <= '0';
            xs(4)  <= '0';
            xs(5)  <= '0';
            xs(6)  <= '1';
            xs(7)  <= '0';
            xs(8)  <= '0';
            xs(9)  <= '0';
            xs(10) <= '0';
            xs(11) <= '0';
            xs(12) <= '0';
            xs(13) <= '0';
            xs(14) <= '0';
            xs(15) <= '0';
            xs(16) <= '0';
            xs(17) <= '0';
            xs(18) <= '0';
            xs(19) <= '0';
            xs(20) <= '0'; 

        when "1000"&"1000" => --t8q8
            xs(0)  <= '0';
            xs(1)  <= '0';
            xs(2)  <= '0';
            xs(3)  <= '0';
            xs(4)  <= '0';
            xs(5)  <= '1';
            xs(6)  <= '0';
            xs(7)  <= '0';
            xs(8)  <= '0';
            xs(9)  <= '0';
            xs(10) <= '0';
            xs(11) <= '0';
            xs(12) <= '0';
            xs(13) <= '0';
            xs(14) <= '0';
            xs(15) <= '0';
            xs(16) <= '0';
            xs(17) <= '0';
            xs(18) <= '0';
            xs(19) <= '0';
            xs(20) <= '0'; 

        when "1000"&"1001" => --t9q8
            xs(0)  <= '0';
            xs(1)  <= '0';
            xs(2)  <= '0';
            xs(3)  <= '0';
            xs(4)  <= '0';
            xs(5)  <= '0';
            xs(6)  <= '0';
            xs(7)  <= '0';
            xs(8)  <= '0';
            xs(9)  <= '0';
            xs(10) <= '0';
            xs(11) <= '0';
            xs(12) <= '0';
            xs(13) <= '0';
            xs(14) <= '1';
            xs(15) <= '0';
            xs(16) <= '0';
            xs(17) <= '0';
            xs(18) <= '0';
            xs(19) <= '0';
            xs(20) <= '0'; 

------------  FIN -> 08h  JMP [DIR]  

------------ 09h  JC DIR   
        --       q & t
        when "1001"&"0000" => --t0
            xs(0)  <= '0';
            xs(1)  <= '0';
            xs(2)  <= '0';
            xs(3)  <= '0';
            xs(4)  <= '0';
            xs(5)  <= '0';
            xs(6)  <= '0';
            xs(7)  <= '0';
            xs(8)  <= '1';
            xs(9)  <= '0';
            xs(10) <= '0';
            xs(11) <= '0';
            xs(12) <= '0';
            xs(13) <= '0';
            xs(14) <= '0';
            xs(15) <= '0';
            xs(16) <= '0';
            xs(17) <= '0';
            xs(18) <= '0';
            xs(19) <= '0';
            xs(20) <= '0';

        when "1001"&"0001" => --t1
            xs(0)  <= '0';
            xs(1)  <= '0';
            xs(2)  <= '1';
            xs(3)  <= '0';
            xs(4)  <= '0';
            xs(5)  <= '0';
            xs(6)  <= '1';
            xs(7)  <= '0';
            xs(8)  <= '0';
            xs(9)  <= '0';
            xs(10) <= '0';
            xs(11) <= '0';
            xs(12) <= '0';
            xs(13) <= '0';
            xs(14) <= '0';
            xs(15) <= '0';
            xs(16) <= '0';
            xs(17) <= '0';
            xs(18) <= '0';
            xs(19) <= '0';
            xs(20) <= '0';    
            
        when "1001"&"0010" => --t2
            xs(0)  <= '1';
            xs(1)  <= '0';
            xs(2)  <= '0';
            xs(3)  <= '0';
            xs(4)  <= '0';
            xs(5)  <= '0';
            xs(6)  <= '0';
            xs(7)  <= '0';
            xs(8)  <= '0';
            xs(9)  <= '0';
            xs(10) <= '0';
            xs(11) <= '0';
            xs(12) <= '0';
            xs(13) <= '0';
            xs(14) <= '0';
            xs(15) <= '0';
            xs(16) <= '0';
            xs(17) <= '0';
            xs(18) <= '0';
            xs(19) <= '0';
            xs(20) <= '0';    
            
        when "1001"&"0011" => --t3q9
            xs(0)  <= '0';
            xs(1)  <= '0';
            xs(2)  <= '0';
            xs(3)  <= '0';
            xs(4)  <= '0';
            xs(5)  <= '0';
            xs(6)  <= '0';
            xs(7)  <= '0';
            xs(8)  <= '1';
            xs(9)  <= '0';
            xs(10) <= '0';
            xs(11) <= '0';
            xs(12) <= '0';
            xs(13) <= '0';
            xs(14) <= '0';
            xs(15) <= '0';
            xs(16) <= '0';
            xs(17) <= '0';
            xs(18) <= '0';
            xs(19) <= '0';
            xs(20) <= '0';  
            
        when "1001"&"0100" => --t4q9
            xs(0)  <= '0';
            xs(1)  <= '0';
            xs(2)  <= '1';
            xs(3)  <= '0';
            xs(4)  <= '0';
            xs(5)  <= '0';
            xs(6)  <= '1';
            xs(7)  <= '0';
            xs(8)  <= '0';
            xs(9)  <= '0';
            xs(10) <= '0';
            xs(11) <= '0';
            xs(12) <= '0';
            xs(13) <= '0';
            xs(14) <= '0';
            xs(15) <= '0';
            xs(16) <= '0';
            xs(17) <= '0';
            xs(18) <= '0';
            xs(19) <= '0';
            xs(20) <= '0';   

        when "1001"&"0101" => --t5q9
            xs(0)  <= '0';
            xs(1)  <= '0';
            xs(2)  <= '0';
            xs(3)  <= '0';
            xs(4)  <= '0';
            xs(5)  <= '0';
            xs(6)  <= '0';
            xs(7)  <= '0';
            xs(8)  <= '0';
            xs(9)  <= '0';
            xs(10) <= '1';
            xs(11) <= '0';
            xs(12) <= '0';
            xs(13) <= '0';
            xs(14) <= '0';
            xs(15) <= '0';
            xs(16) <= '0';
            xs(17) <= '0';
            xs(18) <= '0';
            xs(19) <= '0';
            xs(20) <= '0'; 
            
        when "1001"&"0110" => --t6q9
            xs(0)  <= '0';
            xs(1)  <= '0';
            xs(2)  <= '0';
            xs(3)  <= '0';
            xs(4)  <= '0';
            xs(5)  <= '0';
            xs(6)  <= '0';
            xs(7)  <= '0';
            xs(8)  <= '1';
            xs(9)  <= '0';
            xs(10) <= '0';
            xs(11) <= '0';
            xs(12) <= '0';
            xs(13) <= '0';
            xs(14) <= '0';
            xs(15) <= '0';
            xs(16) <= '0';
            xs(17) <= '0';
            xs(18) <= '0';
            xs(19) <= '0';
            xs(20) <= '0'; 

        when "1001"&"0111" => --t7q9
            xs(0)  <= '0';
            xs(1)  <= '0';
            xs(2)  <= '1';
            xs(3)  <= '0';
            xs(4)  <= '0';
            xs(5)  <= '0';
            xs(6)  <= '1';
            xs(7)  <= '0';
            xs(8)  <= '0';
            xs(9)  <= '0';
            xs(10) <= '0';
            xs(11) <= '0';
            xs(12) <= '0';
            xs(13) <= '0';
            xs(14) <= '0';
            xs(15) <= '0';
            xs(16) <= '0';
            xs(17) <= '0';
            xs(18) <= '0';
            xs(19) <= '0';
            xs(20) <= '0'; 

        when "1001"&"1000" => --t8q9
           if (c_in = '1') then
                xs(0)  <= '0';
                xs(1)  <= '0';
                xs(2)  <= '0';
                xs(3)  <= '0';
                xs(4)  <= '0';
                xs(5)  <= '1';
                xs(6)  <= '0';
                xs(7)  <= '0';
                xs(8)  <= '0';
                xs(9)  <= '0';
                xs(10) <= '0';
                xs(11) <= '0';
                xs(12) <= '0';
                xs(13) <= '0';
                xs(14) <= '0';
                xs(15) <= '0';
                xs(16) <= '0';
                xs(17) <= '0';
                xs(18) <= '0';
                xs(19) <= '0';
                xs(20) <= '0'; 
            else
                xs(0)  <= '0';
                xs(1)  <= '0';
                xs(2)  <= '0';
                xs(3)  <= '0';
                xs(4)  <= '0';
                xs(5)  <= '0';
                xs(6)  <= '0';
                xs(7)  <= '0';
                xs(8)  <= '0';
                xs(9)  <= '0';
                xs(10) <= '0';
                xs(11) <= '0';
                xs(12) <= '0';
                xs(13) <= '0';
                xs(14) <= '1';
                xs(15) <= '0';
                xs(16) <= '0';
                xs(17) <= '0';
                xs(18) <= '0';
                xs(19) <= '0';
                xs(20) <= '0'; 
           end if ;

        when "1001"&"1001" => --t9q9
            xs(0)  <= '0';
            xs(1)  <= '0';
            xs(2)  <= '0';
            xs(3)  <= '0';
            xs(4)  <= '0';
            xs(5)  <= '0';
            xs(6)  <= '0';
            xs(7)  <= '0';
            xs(8)  <= '0';
            xs(9)  <= '0';
            xs(10) <= '0';
            xs(11) <= '0';
            xs(12) <= '0';
            xs(13) <= '0';
            xs(14) <= '1';
            xs(15) <= '0';
            xs(16) <= '0';
            xs(17) <= '0';
            xs(18) <= '0';
            xs(19) <= '0';
            xs(20) <= '0'; 

  
------------  FIN -> 09h  JC DIR    

------------ 0Ah  JZ DIR   
        --       q & t
        when "1010"&"0000" => --t0
            xs(0)  <= '0';
            xs(1)  <= '0';
            xs(2)  <= '0';
            xs(3)  <= '0';
            xs(4)  <= '0';
            xs(5)  <= '0';
            xs(6)  <= '0';
            xs(7)  <= '0';
            xs(8)  <= '1';
            xs(9)  <= '0';
            xs(10) <= '0';
            xs(11) <= '0';
            xs(12) <= '0';
            xs(13) <= '0';
            xs(14) <= '0';
            xs(15) <= '0';
            xs(16) <= '0';
            xs(17) <= '0';
            xs(18) <= '0';
            xs(19) <= '0';
            xs(20) <= '0';

        when "1010"&"0001" => --t1
            xs(0)  <= '0';
            xs(1)  <= '0';
            xs(2)  <= '1';
            xs(3)  <= '0';
            xs(4)  <= '0';
            xs(5)  <= '0';
            xs(6)  <= '1';
            xs(7)  <= '0';
            xs(8)  <= '0';
            xs(9)  <= '0';
            xs(10) <= '0';
            xs(11) <= '0';
            xs(12) <= '0';
            xs(13) <= '0';
            xs(14) <= '0';
            xs(15) <= '0';
            xs(16) <= '0';
            xs(17) <= '0';
            xs(18) <= '0';
            xs(19) <= '0';
            xs(20) <= '0';    
            
        when "1010"&"0010" => --t2
            xs(0)  <= '1';
            xs(1)  <= '0';
            xs(2)  <= '0';
            xs(3)  <= '0';
            xs(4)  <= '0';
            xs(5)  <= '0';
            xs(6)  <= '0';
            xs(7)  <= '0';
            xs(8)  <= '0';
            xs(9)  <= '0';
            xs(10) <= '0';
            xs(11) <= '0';
            xs(12) <= '0';
            xs(13) <= '0';
            xs(14) <= '0';
            xs(15) <= '0';
            xs(16) <= '0';
            xs(17) <= '0';
            xs(18) <= '0';
            xs(19) <= '0';
            xs(20) <= '0';    
            
        when "1010"&"0011" => --t3qA
            xs(0)  <= '0';
            xs(1)  <= '0';
            xs(2)  <= '0';
            xs(3)  <= '0';
            xs(4)  <= '0';
            xs(5)  <= '0';
            xs(6)  <= '0';
            xs(7)  <= '0';
            xs(8)  <= '1';
            xs(9)  <= '0';
            xs(10) <= '0';
            xs(11) <= '0';
            xs(12) <= '0';
            xs(13) <= '0';
            xs(14) <= '0';
            xs(15) <= '0';
            xs(16) <= '0';
            xs(17) <= '0';
            xs(18) <= '0';
            xs(19) <= '0';
            xs(20) <= '0';  
            
        when "1010"&"0100" => --t4qA
            xs(0)  <= '0';
            xs(1)  <= '0';
            xs(2)  <= '1';
            xs(3)  <= '0';
            xs(4)  <= '0';
            xs(5)  <= '0';
            xs(6)  <= '1';
            xs(7)  <= '0';
            xs(8)  <= '0';
            xs(9)  <= '0';
            xs(10) <= '0';
            xs(11) <= '0';
            xs(12) <= '0';
            xs(13) <= '0';
            xs(14) <= '0';
            xs(15) <= '0';
            xs(16) <= '0';
            xs(17) <= '0';
            xs(18) <= '0';
            xs(19) <= '0';
            xs(20) <= '0';   

        when "1010"&"0101" => --t5qA
            xs(0)  <= '0';
            xs(1)  <= '0';
            xs(2)  <= '0';
            xs(3)  <= '0';
            xs(4)  <= '0';
            xs(5)  <= '0';
            xs(6)  <= '0';
            xs(7)  <= '0';
            xs(8)  <= '0';
            xs(9)  <= '0';
            xs(10) <= '1';
            xs(11) <= '0';
            xs(12) <= '0';
            xs(13) <= '0';
            xs(14) <= '0';
            xs(15) <= '0';
            xs(16) <= '0';
            xs(17) <= '0';
            xs(18) <= '0';
            xs(19) <= '0';
            xs(20) <= '0'; 
            
        when "1010"&"0110" => --t6qA
            xs(0)  <= '0';
            xs(1)  <= '0';
            xs(2)  <= '0';
            xs(3)  <= '0';
            xs(4)  <= '0';
            xs(5)  <= '0';
            xs(6)  <= '0';
            xs(7)  <= '0';
            xs(8)  <= '1';
            xs(9)  <= '0';
            xs(10) <= '0';
            xs(11) <= '0';
            xs(12) <= '0';
            xs(13) <= '0';
            xs(14) <= '0';
            xs(15) <= '0';
            xs(16) <= '0';
            xs(17) <= '0';
            xs(18) <= '0';
            xs(19) <= '0';
            xs(20) <= '0'; 

        when "1010"&"0111" => --t7qA
            xs(0)  <= '0';
            xs(1)  <= '0';
            xs(2)  <= '1';
            xs(3)  <= '0';
            xs(4)  <= '0';
            xs(5)  <= '0';
            xs(6)  <= '1';
            xs(7)  <= '0';
            xs(8)  <= '0';
            xs(9)  <= '0';
            xs(10) <= '0';
            xs(11) <= '0';
            xs(12) <= '0';
            xs(13) <= '0';
            xs(14) <= '0';
            xs(15) <= '0';
            xs(16) <= '0';
            xs(17) <= '0';
            xs(18) <= '0';
            xs(19) <= '0';
            xs(20) <= '0'; 

        when "1010"&"1000" => --t8qA
           if (z_in = '1') then
                xs(0)  <= '0';
                xs(1)  <= '0';
                xs(2)  <= '0';
                xs(3)  <= '0';
                xs(4)  <= '0';
                xs(5)  <= '1';
                xs(6)  <= '0';
                xs(7)  <= '0';
                xs(8)  <= '0';
                xs(9)  <= '0';
                xs(10) <= '0';
                xs(11) <= '0';
                xs(12) <= '0';
                xs(13) <= '0';
                xs(14) <= '0';
                xs(15) <= '0';
                xs(16) <= '0';
                xs(17) <= '0';
                xs(18) <= '0';
                xs(19) <= '0';
                xs(20) <= '0'; 
            else
                xs(0)  <= '0';
                xs(1)  <= '0';
                xs(2)  <= '0';
                xs(3)  <= '0';
                xs(4)  <= '0';
                xs(5)  <= '0';
                xs(6)  <= '0';
                xs(7)  <= '0';
                xs(8)  <= '0';
                xs(9)  <= '0';
                xs(10) <= '0';
                xs(11) <= '0';
                xs(12) <= '0';
                xs(13) <= '0';
                xs(14) <= '1';
                xs(15) <= '0';
                xs(16) <= '0';
                xs(17) <= '0';
                xs(18) <= '0';
                xs(19) <= '0';
                xs(20) <= '0'; 
           end if ;

        when "1010"&"1001" => --t9qA
            xs(0)  <= '0';
            xs(1)  <= '0';
            xs(2)  <= '0';
            xs(3)  <= '0';
            xs(4)  <= '0';
            xs(5)  <= '0';
            xs(6)  <= '0';
            xs(7)  <= '0';
            xs(8)  <= '0';
            xs(9)  <= '0';
            xs(10) <= '0';
            xs(11) <= '0';
            xs(12) <= '0';
            xs(13) <= '0';
            xs(14) <= '1';
            xs(15) <= '0';
            xs(16) <= '0';
            xs(17) <= '0';
            xs(18) <= '0';
            xs(19) <= '0';
            xs(20) <= '0'; 

  
------------  FIN -> 0Ah  JZ DIR  

------------ 0Bh  JSR DIR   
        --       q & t
        when "1011"&"0000" => --t0
            xs(0)  <= '0';
            xs(1)  <= '0';
            xs(2)  <= '0';
            xs(3)  <= '0';
            xs(4)  <= '0';
            xs(5)  <= '0';
            xs(6)  <= '0';
            xs(7)  <= '0';
            xs(8)  <= '1';
            xs(9)  <= '0';
            xs(10) <= '0';
            xs(11) <= '0';
            xs(12) <= '0';
            xs(13) <= '0';
            xs(14) <= '0';
            xs(15) <= '0';
            xs(16) <= '0';
            xs(17) <= '0';
            xs(18) <= '0';
            xs(19) <= '0';
            xs(20) <= '0';

        when "1011"&"0001" => --t1
            xs(0)  <= '0';
            xs(1)  <= '0';
            xs(2)  <= '1';
            xs(3)  <= '0';
            xs(4)  <= '0';
            xs(5)  <= '0';
            xs(6)  <= '1';
            xs(7)  <= '0';
            xs(8)  <= '0';
            xs(9)  <= '0';
            xs(10) <= '0';
            xs(11) <= '0';
            xs(12) <= '0';
            xs(13) <= '0';
            xs(14) <= '0';
            xs(15) <= '0';
            xs(16) <= '0';
            xs(17) <= '0';
            xs(18) <= '0';
            xs(19) <= '0';
            xs(20) <= '0';    
            
        when "1011"&"0010" => --t2
            xs(0)  <= '1';
            xs(1)  <= '0';
            xs(2)  <= '0';
            xs(3)  <= '0';
            xs(4)  <= '0';
            xs(5)  <= '0';
            xs(6)  <= '0';
            xs(7)  <= '0';
            xs(8)  <= '0';
            xs(9)  <= '0';
            xs(10) <= '0';
            xs(11) <= '0';
            xs(12) <= '0';
            xs(13) <= '0';
            xs(14) <= '0';
            xs(15) <= '0';
            xs(16) <= '0';
            xs(17) <= '0';
            xs(18) <= '0';
            xs(19) <= '0';
            xs(20) <= '0';    
            
        when "1011"&"0011" => --t3qB
            xs(0)  <= '0';
            xs(1)  <= '0';
            xs(2)  <= '0';
            xs(3)  <= '0';
            xs(4)  <= '0';
            xs(5)  <= '0';
            xs(6)  <= '0';
            xs(7)  <= '0';
            xs(8)  <= '1';
            xs(9)  <= '0';
            xs(10) <= '0';
            xs(11) <= '0';
            xs(12) <= '0';
            xs(13) <= '0';
            xs(14) <= '0';
            xs(15) <= '0';
            xs(16) <= '0';
            xs(17) <= '0';
            xs(18) <= '0';
            xs(19) <= '0';
            xs(20) <= '0';  
            
        when "1011"&"0100" => --t4qB
            xs(0)  <= '0';
            xs(1)  <= '0';
            xs(2)  <= '1';
            xs(3)  <= '0';
            xs(4)  <= '0';
            xs(5)  <= '0';
            xs(6)  <= '1';
            xs(7)  <= '0';
            xs(8)  <= '0';
            xs(9)  <= '0';
            xs(10) <= '0';
            xs(11) <= '0';
            xs(12) <= '0';
            xs(13) <= '0';
            xs(14) <= '0';
            xs(15) <= '0';
            xs(16) <= '0';
            xs(17) <= '0';
            xs(18) <= '0';
            xs(19) <= '0';
            xs(20) <= '0';   

        when "1011"&"0101" => --t5qB
            xs(0)  <= '0';
            xs(1)  <= '0';
            xs(2)  <= '0';
            xs(3)  <= '0';
            xs(4)  <= '0';
            xs(5)  <= '0';
            xs(6)  <= '0';
            xs(7)  <= '0';
            xs(8)  <= '1';
            xs(9)  <= '0';
            xs(10) <= '1';
            xs(11) <= '0';
            xs(12) <= '0';
            xs(13) <= '0';
            xs(14) <= '0';
            xs(15) <= '0';
            xs(16) <= '0';
            xs(17) <= '0';
            xs(18) <= '0';
            xs(19) <= '0';
            xs(20) <= '0'; 
            
        when "1011"&"0110" => --t6qB
            xs(0)  <= '0';
            xs(1)  <= '0';
            xs(2)  <= '1';
            xs(3)  <= '0';
            xs(4)  <= '0';
            xs(5)  <= '0';
            xs(6)  <= '1';
            xs(7)  <= '0';
            xs(8)  <= '0';
            xs(9)  <= '0';
            xs(10) <= '0';
            xs(11) <= '0';
            xs(12) <= '0';
            xs(13) <= '0';
            xs(14) <= '0';
            xs(15) <= '0';
            xs(16) <= '0';
            xs(17) <= '0';
            xs(18) <= '0';
            xs(19) <= '0';
            xs(20) <= '0'; 

        when "1011"&"0111" => --t7qB
            xs(0)  <= '0';
            xs(1)  <= '0';
            xs(2)  <= '0';
            xs(3)  <= '0';
            xs(4)  <= '0';
            xs(5)  <= '0';
            xs(6)  <= '0';
            xs(7)  <= '0';
            xs(8)  <= '0';
            xs(9)  <= '1';
            xs(10) <= '0';
            xs(11) <= '0';
            xs(12) <= '0';
            xs(13) <= '0';
            xs(14) <= '0';
            xs(15) <= '1';
            xs(16) <= '1';
            xs(17) <= '1';
            xs(18) <= '0';
            xs(19) <= '1';
            xs(20) <= '0'; 

        when "1011"&"1000" => --t8qB
                xs(0)  <= '0';
                xs(1)  <= '0';
                xs(2)  <= '0';
                xs(3)  <= '1';
                xs(4)  <= '0';
                xs(5)  <= '0';
                xs(6)  <= '0';
                xs(7)  <= '0';
                xs(8)  <= '0';
                xs(9)  <= '0';
                xs(10) <= '0';
                xs(11) <= '0';
                xs(12) <= '0';
                xs(13) <= '1';
                xs(14) <= '0';
                xs(15) <= '0';
                xs(16) <= '0';
                xs(17) <= '0';
                xs(18) <= '0';
                xs(19) <= '0';
                xs(20) <= '0'; 

        when "1011"&"1001" => --t9qB
            xs(0)  <= '0';
            xs(1)  <= '0';
            xs(2)  <= '0';
            xs(3)  <= '0';
            xs(4)  <= '0';
            xs(5)  <= '0';
            xs(6)  <= '0';
            xs(7)  <= '0';
            xs(8)  <= '0';
            xs(9)  <= '0';
            xs(10) <= '0';
            xs(11) <= '0';
            xs(12) <= '0';
            xs(13) <= '0';
            xs(14) <= '0';
            xs(15) <= '0';
            xs(16) <= '0';
            xs(17) <= '0';
            xs(18) <= '0';
            xs(19) <= '0';
            xs(20) <= '1'; 

        when "1011"&"1010" => --tAqB
            xs(0)  <= '0';
            xs(1)  <= '0';
            xs(2)  <= '0';
            xs(3)  <= '0';
            xs(4)  <= '0';
            xs(5)  <= '0';
            xs(6)  <= '0';
            xs(7)  <= '0';
            xs(8)  <= '0';
            xs(9)  <= '1';
            xs(10) <= '0';
            xs(11) <= '0';
            xs(12) <= '0';
            xs(13) <= '0';
            xs(14) <= '0';
            xs(15) <= '0';
            xs(16) <= '0';
            xs(17) <= '0';
            xs(18) <= '0';
            xs(19) <= '0';
            xs(20) <= '0'; 
  
        when "1011"&"1011" => --tBqB
            xs(0)  <= '0';
            xs(1)  <= '0';
            xs(2)  <= '0';
            xs(3)  <= '0';
            xs(4)  <= '1';
            xs(5)  <= '0';
            xs(6)  <= '0';
            xs(7)  <= '0';
            xs(8)  <= '0';
            xs(9)  <= '0';
            xs(10) <= '0';
            xs(11) <= '0';
            xs(12) <= '0';
            xs(13) <= '1';
            xs(14) <= '0';
            xs(15) <= '0';
            xs(16) <= '0';
            xs(17) <= '0';
            xs(18) <= '0';
            xs(19) <= '0';
            xs(20) <= '0';
            
        when "1011"&"1100" => --tCqB
            xs(0)  <= '0';
            xs(1)  <= '0';
            xs(2)  <= '0';
            xs(3)  <= '0';
            xs(4)  <= '0';
            xs(5)  <= '0';
            xs(6)  <= '0';
            xs(7)  <= '0';
            xs(8)  <= '0';
            xs(9)  <= '0';
            xs(10) <= '0';
            xs(11) <= '0';
            xs(12) <= '0';
            xs(13) <= '0';
            xs(14) <= '0';
            xs(15) <= '0';
            xs(16) <= '0';
            xs(17) <= '0';
            xs(18) <= '0';
            xs(19) <= '0';
            xs(20) <= '1';
            
        when "1011"&"1101" => --tDqB
            xs(0)  <= '0';
            xs(1)  <= '1';
            xs(2)  <= '0';
            xs(3)  <= '0';
            xs(4)  <= '0';
            xs(5)  <= '0';
            xs(6)  <= '0';
            xs(7)  <= '0';
            xs(8)  <= '0';
            xs(9)  <= '0';
            xs(10) <= '0';
            xs(11) <= '0';
            xs(12) <= '0';
            xs(13) <= '0';
            xs(14) <= '0';
            xs(15) <= '0';
            xs(16) <= '0';
            xs(17) <= '0';
            xs(18) <= '0';
            xs(19) <= '0';
            xs(20) <= '0'; 

        when "1011"&"1110" => --tEqB
            xs(0)  <= '0';
            xs(1)  <= '0';
            xs(2)  <= '0';
            xs(3)  <= '0';
            xs(4)  <= '0';
            xs(5)  <= '1';
            xs(6)  <= '0';
            xs(7)  <= '0';
            xs(8)  <= '0';
            xs(9)  <= '0';
            xs(10) <= '0';
            xs(11) <= '0';
            xs(12) <= '0';
            xs(13) <= '0';
            xs(14) <= '0';
            xs(15) <= '0';
            xs(16) <= '0';
            xs(17) <= '0';
            xs(18) <= '0';
            xs(19) <= '0';
            xs(20) <= '0'; 

        when "1011"&"1111" => --tFqB
            xs(0)  <= '0';
            xs(1)  <= '0';
            xs(2)  <= '0';
            xs(3)  <= '0';
            xs(4)  <= '0';
            xs(5)  <= '0';
            xs(6)  <= '0';
            xs(7)  <= '0';
            xs(8)  <= '0';
            xs(9)  <= '0';
            xs(10) <= '0';
            xs(11) <= '0';
            xs(12) <= '0';
            xs(13) <= '0';
            xs(14) <= '1';
            xs(15) <= '0';
            xs(16) <= '0';
            xs(17) <= '0';
            xs(18) <= '0';
            xs(19) <= '0';
            xs(20) <= '0'; 
------------  FIN -> 0Bh  JSR DIR  

------------ 0Ch  RTS 
        --       q & t
        when "1100"&"00000" => --t0
            xs(0)  <= '0';
            xs(1)  <= '0';
            xs(2)  <= '0';
            xs(3)  <= '0';
            xs(4)  <= '0';
            xs(5)  <= '0';
            xs(6)  <= '0';
            xs(7)  <= '0';
            xs(8)  <= '1';
            xs(9)  <= '0';
            xs(10) <= '0';
            xs(11) <= '0';
            xs(12) <= '0';
            xs(13) <= '0';
            xs(14) <= '0';
            xs(15) <= '0';
            xs(16) <= '0';
            xs(17) <= '0';
            xs(18) <= '0';
            xs(19) <= '0';
            xs(20) <= '0';

        when "1100"&"00001" => --t1
            xs(0)  <= '0';
            xs(1)  <= '0';
            xs(2)  <= '1';
            xs(3)  <= '0';
            xs(4)  <= '0';
            xs(5)  <= '0';
            xs(6)  <= '1';
            xs(7)  <= '0';
            xs(8)  <= '0';
            xs(9)  <= '0';
            xs(10) <= '0';
            xs(11) <= '0';
            xs(12) <= '0';
            xs(13) <= '0';
            xs(14) <= '0';
            xs(15) <= '0';
            xs(16) <= '0';
            xs(17) <= '0';
            xs(18) <= '0';
            xs(19) <= '0';
            xs(20) <= '0';    
            
        when "1100"&"00010" => --t2
            xs(0)  <= '1';
            xs(1)  <= '0';
            xs(2)  <= '0';
            xs(3)  <= '0';
            xs(4)  <= '0';
            xs(5)  <= '0';
            xs(6)  <= '0';
            xs(7)  <= '0';
            xs(8)  <= '0';
            xs(9)  <= '0';
            xs(10) <= '0';
            xs(11) <= '0';
            xs(12) <= '0';
            xs(13) <= '0';
            xs(14) <= '0';
            xs(15) <= '0';
            xs(16) <= '0';
            xs(17) <= '0';
            xs(18) <= '0';
            xs(19) <= '0';
            xs(20) <= '0';    
            
        when "1100"&"00011" => --t3qC
            xs(0)  <= '0';
            xs(1)  <= '0';
            xs(2)  <= '0';
            xs(3)  <= '0';
            xs(4)  <= '0';
            xs(5)  <= '0';
            xs(6)  <= '0';
            xs(7)  <= '0';
            xs(8)  <= '0';
            xs(9)  <= '0';
            xs(10) <= '0';
            xs(11) <= '0';
            xs(12) <= '1';
            xs(13) <= '0';
            xs(14) <= '0';
            xs(15) <= '0';
            xs(16) <= '0';
            xs(17) <= '0';
            xs(18) <= '0';
            xs(19) <= '0';
            xs(20) <= '0';  
            
        when "1100"&"00100" => --t4qC
            xs(0)  <= '0';
            xs(1)  <= '0';
            xs(2)  <= '0';
            xs(3)  <= '0';
            xs(4)  <= '0';
            xs(5)  <= '0';
            xs(6)  <= '0';
            xs(7)  <= '0';
            xs(8)  <= '0';
            xs(9)  <= '1';
            xs(10) <= '0';
            xs(11) <= '0';
            xs(12) <= '0';
            xs(13) <= '0';
            xs(14) <= '0';
            xs(15) <= '0';
            xs(16) <= '0';
            xs(17) <= '0';
            xs(18) <= '0';
            xs(19) <= '0';
            xs(20) <= '0';   

        when "1100"&"00101" => --t5qC
            xs(0)  <= '0';
            xs(1)  <= '0';
            xs(2)  <= '1';
            xs(3)  <= '0';
            xs(4)  <= '0';
            xs(5)  <= '0';
            xs(6)  <= '0';
            xs(7)  <= '0';
            xs(8)  <= '1';
            xs(9)  <= '0';
            xs(10) <= '0';
            xs(11) <= '0';
            xs(12) <= '1';
            xs(13) <= '0';
            xs(14) <= '0';
            xs(15) <= '0';
            xs(16) <= '0';
            xs(17) <= '0';
            xs(18) <= '0';
            xs(19) <= '0';
            xs(20) <= '0'; 
            
        when "1100"&"00110" => --t6qC
            xs(0)  <= '0';
            xs(1)  <= '0';
            xs(2)  <= '0';
            xs(3)  <= '0';
            xs(4)  <= '0';
            xs(5)  <= '0';
            xs(6)  <= '0';
            xs(7)  <= '0';
            xs(8)  <= '0';
            xs(9)  <= '0';
            xs(10) <= '1';
            xs(11) <= '0';
            xs(12) <= '0';
            xs(13) <= '0';
            xs(14) <= '0';
            xs(15) <= '0';
            xs(16) <= '0';
            xs(17) <= '0';
            xs(18) <= '0';
            xs(19) <= '0';
            xs(20) <= '0'; 

        when "1100"&"00110" => --t7qC
            xs(0)  <= '0';
            xs(1)  <= '0';
            xs(2)  <= '0';
            xs(3)  <= '0';
            xs(4)  <= '0';
            xs(5)  <= '0';
            xs(6)  <= '0';
            xs(7)  <= '0';
            xs(8)  <= '0';
            xs(9)  <= '1';
            xs(10) <= '0';
            xs(11) <= '0';
            xs(12) <= '0';
            xs(13) <= '0';
            xs(14) <= '0';
            xs(15) <= '0';
            xs(16) <= '0';
            xs(17) <= '0';
            xs(18) <= '0';
            xs(19) <= '0';
            xs(20) <= '0'; 

        when "1100"&"00111" => --t8qC
                xs(0)  <= '0';
                xs(1)  <= '0';
                xs(2)  <= '1';
                xs(3)  <= '0';
                xs(4)  <= '0';
                xs(5)  <= '0';
                xs(6)  <= '0';
                xs(7)  <= '0';
                xs(8)  <= '0';
                xs(9)  <= '1';
                xs(10) <= '0';
                xs(11) <= '0';
                xs(12) <= '0';
                xs(13) <= '0';
                xs(14) <= '0';
                xs(15) <= '0';
                xs(16) <= '0';
                xs(17) <= '0';
                xs(18) <= '0';
                xs(19) <= '0';
                xs(20) <= '0'; 

        when "1100"&"01000" => --t9qC
            xs(0)  <= '0';
            xs(1)  <= '0';
            xs(2)  <= '0';
            xs(3)  <= '0';
            xs(4)  <= '0';
            xs(5)  <= '1';
            xs(6)  <= '0';
            xs(7)  <= '0';
            xs(8)  <= '0';
            xs(9)  <= '0';
            xs(10) <= '0';
            xs(11) <= '0';
            xs(12) <= '0';
            xs(13) <= '0';
            xs(14) <= '0';
            xs(15) <= '0';
            xs(16) <= '0';
            xs(17) <= '0';
            xs(18) <= '0';
            xs(19) <= '0';
            xs(20) <= '0'; 

        when "1100"&"01001" => --tAqC
            xs(0)  <= '0';
            xs(1)  <= '0';
            xs(2)  <= '0';
            xs(3)  <= '0';
            xs(4)  <= '0';
            xs(5)  <= '0';
            xs(6)  <= '0';
            xs(7)  <= '0';
            xs(8)  <= '0';
            xs(9)  <= '0';
            xs(10) <= '0';
            xs(11) <= '0';
            xs(12) <= '0';
            xs(13) <= '0';
            xs(14) <= '1';
            xs(15) <= '0';
            xs(16) <= '0';
            xs(17) <= '0';
            xs(18) <= '0';
            xs(19) <= '0';
            xs(20) <= '0'; 
------------  FIN -> 0Ch  RTS  

------------  0Dh  LSL A 
        --       q & t
        when "1100"&"0000" => --t0
            xs(0)  <= '0';
            xs(1)  <= '0';
            xs(2)  <= '0';
            xs(3)  <= '0';
            xs(4)  <= '0';
            xs(5)  <= '0';
            xs(6)  <= '0';
            xs(7)  <= '0';
            xs(8)  <= '1';
            xs(9)  <= '0';
            xs(10) <= '0';
            xs(11) <= '0';
            xs(12) <= '0';
            xs(13) <= '0';
            xs(14) <= '0';
            xs(15) <= '0';
            xs(16) <= '0';
            xs(17) <= '0';
            xs(18) <= '0';
            xs(19) <= '0';
            xs(20) <= '0';

        when "1100"&"0001" => --t1
            xs(0)  <= '0';
            xs(1)  <= '0';
            xs(2)  <= '1';
            xs(3)  <= '0';
            xs(4)  <= '0';
            xs(5)  <= '0';
            xs(6)  <= '1';
            xs(7)  <= '0';
            xs(8)  <= '0';
            xs(9)  <= '0';
            xs(10) <= '0';
            xs(11) <= '0';
            xs(12) <= '0';
            xs(13) <= '0';
            xs(14) <= '0';
            xs(15) <= '0';
            xs(16) <= '0';
            xs(17) <= '0';
            xs(18) <= '0';
            xs(19) <= '0';
            xs(20) <= '0';    
            
        when "1100"&"0010" => --t2
            xs(0)  <= '1';
            xs(1)  <= '0';
            xs(2)  <= '0';
            xs(3)  <= '0';
            xs(4)  <= '0';
            xs(5)  <= '0';
            xs(6)  <= '0';
            xs(7)  <= '0';
            xs(8)  <= '0';
            xs(9)  <= '0';
            xs(10) <= '0';
            xs(11) <= '0';
            xs(12) <= '0';
            xs(13) <= '0';
            xs(14) <= '0';
            xs(15) <= '0';
            xs(16) <= '0';
            xs(17) <= '0';
            xs(18) <= '0';
            xs(19) <= '0';
            xs(20) <= '0';    
            
        when "1100"&"0011" => --t3qD
            xs(0)  <= '0';
            xs(1)  <= '0';
            xs(2)  <= '0';
            xs(3)  <= '0';
            xs(4)  <= '0';
            xs(5)  <= '0';
            xs(6)  <= '0';
            xs(7)  <= '0';
            xs(8)  <= '0';
            xs(9)  <= '0';
            xs(10) <= '0';
            xs(11) <= '0';
            xs(12) <= '0';
            xs(13) <= '0';
            xs(14) <= '0';
            xs(15) <= '0';
            xs(16) <= '0';
            xs(17) <= '1';
            xs(18) <= '0';
            xs(19) <= '1';
            xs(20) <= '0';  
            
        when "1100"&"0100" => --t4qD
            xs(0)  <= '0';
            xs(1)  <= '0';
            xs(2)  <= '0';
            xs(3)  <= '0';
            xs(4)  <= '0';
            xs(5)  <= '0';
            xs(6)  <= '0';
            xs(7)  <= '0';
            xs(8)  <= '0';
            xs(9)  <= '0';
            xs(10) <= '0';
            xs(11) <= '0';
            xs(12) <= '0';
            xs(13) <= '0';
            xs(14) <= '1';
            xs(15) <= '0';
            xs(16) <= '0';
            xs(17) <= '0';
            xs(18) <= '0';
            xs(19) <= '0';
            xs(20) <= '0';   
------------  FIN -> 0Dh  LSL A  


------------  0Eh  LSR A 
        --       q & t
        when "1110"&"0000" => --t0
            xs(0)  <= '0';
            xs(1)  <= '0';
            xs(2)  <= '0';
            xs(3)  <= '0';
            xs(4)  <= '0';
            xs(5)  <= '0';
            xs(6)  <= '0';
            xs(7)  <= '0';
            xs(8)  <= '1';
            xs(9)  <= '0';
            xs(10) <= '0';
            xs(11) <= '0';
            xs(12) <= '0';
            xs(13) <= '0';
            xs(14) <= '0';
            xs(15) <= '0';
            xs(16) <= '0';
            xs(17) <= '0';
            xs(18) <= '0';
            xs(19) <= '0';
            xs(20) <= '0';

        when "1110"&"0001" => --t1
            xs(0)  <= '0';
            xs(1)  <= '0';
            xs(2)  <= '1';
            xs(3)  <= '0';
            xs(4)  <= '0';
            xs(5)  <= '0';
            xs(6)  <= '1';
            xs(7)  <= '0';
            xs(8)  <= '0';
            xs(9)  <= '0';
            xs(10) <= '0';
            xs(11) <= '0';
            xs(12) <= '0';
            xs(13) <= '0';
            xs(14) <= '0';
            xs(15) <= '0';
            xs(16) <= '0';
            xs(17) <= '0';
            xs(18) <= '0';
            xs(19) <= '0';
            xs(20) <= '0';    
            
        when "1110"&"0010" => --t2
            xs(0)  <= '1';
            xs(1)  <= '0';
            xs(2)  <= '0';
            xs(3)  <= '0';
            xs(4)  <= '0';
            xs(5)  <= '0';
            xs(6)  <= '0';
            xs(7)  <= '0';
            xs(8)  <= '0';
            xs(9)  <= '0';
            xs(10) <= '0';
            xs(11) <= '0';
            xs(12) <= '0';
            xs(13) <= '0';
            xs(14) <= '0';
            xs(15) <= '0';
            xs(16) <= '0';
            xs(17) <= '0';
            xs(18) <= '0';
            xs(19) <= '0';
            xs(20) <= '0';    
            
        when "1110"&"0011" => --t3qE
            xs(0)  <= '0';
            xs(1)  <= '0';
            xs(2)  <= '0';
            xs(3)  <= '0';
            xs(4)  <= '0';
            xs(5)  <= '0';
            xs(6)  <= '0';
            xs(7)  <= '0';
            xs(8)  <= '0';
            xs(9)  <= '0';
            xs(10) <= '0';
            xs(11) <= '0';
            xs(12) <= '0';
            xs(13) <= '0';
            xs(14) <= '0';
            xs(15) <= '1';
            xs(16) <= '0';
            xs(17) <= '1';
            xs(18) <= '0';
            xs(19) <= '1';
            xs(20) <= '0';  
            
        when "1110"&"0100" => --t4qE
            xs(0)  <= '0';
            xs(1)  <= '0';
            xs(2)  <= '0';
            xs(3)  <= '0';
            xs(4)  <= '0';
            xs(5)  <= '0';
            xs(6)  <= '0';
            xs(7)  <= '0';
            xs(8)  <= '0';
            xs(9)  <= '0';
            xs(10) <= '0';
            xs(11) <= '0';
            xs(12) <= '0';
            xs(13) <= '0';
            xs(14) <= '1';
            xs(15) <= '0';
            xs(16) <= '0';
            xs(17) <= '0';
            xs(18) <= '0';
            xs(19) <= '0';
            xs(20) <= '0';   
------------  FIN -> 0Eh  LSR A  

------------  0Eh  NOT A 
        --       q & t
        when "1111"&"0000" => --t0
            xs(0)  <= '0';
            xs(1)  <= '0';
            xs(2)  <= '0';
            xs(3)  <= '0';
            xs(4)  <= '0';
            xs(5)  <= '0';
            xs(6)  <= '0';
            xs(7)  <= '0';
            xs(8)  <= '1';
            xs(9)  <= '0';
            xs(10) <= '0';
            xs(11) <= '0';
            xs(12) <= '0';
            xs(13) <= '0';
            xs(14) <= '0';
            xs(15) <= '0';
            xs(16) <= '0';
            xs(17) <= '0';
            xs(18) <= '0';
            xs(19) <= '0';
            xs(20) <= '0';

        when "1111"&"0001" => --t1
            xs(0)  <= '0';
            xs(1)  <= '0';
            xs(2)  <= '1';
            xs(3)  <= '0';
            xs(4)  <= '0';
            xs(5)  <= '0';
            xs(6)  <= '1';
            xs(7)  <= '0';
            xs(8)  <= '0';
            xs(9)  <= '0';
            xs(10) <= '0';
            xs(11) <= '0';
            xs(12) <= '0';
            xs(13) <= '0';
            xs(14) <= '0';
            xs(15) <= '0';
            xs(16) <= '0';
            xs(17) <= '0';
            xs(18) <= '0';
            xs(19) <= '0';
            xs(20) <= '0';    
            
        when "1111"&"0010" => --t2
            xs(0)  <= '1';
            xs(1)  <= '0';
            xs(2)  <= '0';
            xs(3)  <= '0';
            xs(4)  <= '0';
            xs(5)  <= '0';
            xs(6)  <= '0';
            xs(7)  <= '0';
            xs(8)  <= '0';
            xs(9)  <= '0';
            xs(10) <= '0';
            xs(11) <= '0';
            xs(12) <= '0';
            xs(13) <= '0';
            xs(14) <= '0';
            xs(15) <= '0';
            xs(16) <= '0';
            xs(17) <= '0';
            xs(18) <= '0';
            xs(19) <= '0';
            xs(20) <= '0';    
            
        when "1111"&"0011" => --t3qF
            xs(0)  <= '0';
            xs(1)  <= '0';
            xs(2)  <= '0';
            xs(3)  <= '0';
            xs(4)  <= '0';
            xs(5)  <= '0';
            xs(6)  <= '0';
            xs(7)  <= '0';
            xs(8)  <= '0';
            xs(9)  <= '0';
            xs(10) <= '0';
            xs(11) <= '0';
            xs(12) <= '0';
            xs(13) <= '0';
            xs(14) <= '0';
            xs(15) <= '0';
            xs(16) <= '0';
            xs(17) <= '1';
            xs(18) <= '0';
            xs(19) <= '1';
            xs(20) <= '0';  
            
        when "1111"&"0100" => --t4qF
            xs(0)  <= '0';
            xs(1)  <= '0';
            xs(2)  <= '0';
            xs(3)  <= '0';
            xs(4)  <= '0';
            xs(5)  <= '0';
            xs(6)  <= '0';
            xs(7)  <= '0';
            xs(8)  <= '0';
            xs(9)  <= '0';
            xs(10) <= '0';
            xs(11) <= '0';
            xs(12) <= '0';
            xs(13) <= '0';
            xs(14) <= '1';
            xs(15) <= '0';
            xs(16) <= '0';
            xs(17) <= '0';
            xs(18) <= '0';
            xs(19) <= '0';
            xs(20) <= '0';   
------------  FIN -> 0Fh  NOT A  
when others =>
        xs <= (others => '0'); --RESET
        end case ;
           
    end process;
   Xs_out <= xs     
end architecture ;


